netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:age.enabled = "no";
    pism_overrides:age.enabled_doc = "Solve age equation (advection equation for ice age).";
    pism_overrides:age.enabled_option = "age";
    pism_overrides:age.enabled_type = "flag";

    pism_overrides:age.initial_value = 0.0;
    pism_overrides:age.initial_value_doc = "Initial age of ice";
    pism_overrides:age.initial_value_type = "number";
    pism_overrides:age.initial_value_units = "years";

    pism_overrides:atmosphere.anomaly.file = "";
    pism_overrides:atmosphere.anomaly.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:atmosphere.anomaly.file_option = "atmosphere_anomaly_file";
    pism_overrides:atmosphere.anomaly.file_type = "string";

    pism_overrides:atmosphere.anomaly.period = 0;
    pism_overrides:atmosphere.anomaly.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.anomaly.period_option = "atmosphere_anomaly_period";
    pism_overrides:atmosphere.anomaly.period_type = "integer";
    pism_overrides:atmosphere.anomaly.period_units = "years";

    pism_overrides:atmosphere.anomaly.reference_year = 0;
    pism_overrides:atmosphere.anomaly.reference_year_doc = "Reference year to use when ``atmosphere.anomaly.period`` is active.";
    pism_overrides:atmosphere.anomaly.reference_year_option = "atmosphere_anomaly_reference_year";
    pism_overrides:atmosphere.anomaly.reference_year_type = "integer";
    pism_overrides:atmosphere.anomaly.reference_year_units = "years";

    pism_overrides:atmosphere.delta_P.file = "";
    pism_overrides:atmosphere.delta_P.file_doc = "Name of the file containing scalar precipitation offsets.";
    pism_overrides:atmosphere.delta_P.file_option = "atmosphere_delta_P_file";
    pism_overrides:atmosphere.delta_P.file_type = "string";

    pism_overrides:atmosphere.delta_P.period = 0;
    pism_overrides:atmosphere.delta_P.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.delta_P.period_option = "atmosphere_delta_P_period";
    pism_overrides:atmosphere.delta_P.period_type = "integer";
    pism_overrides:atmosphere.delta_P.period_units = "years";

    pism_overrides:atmosphere.delta_P.reference_year = 0;
    pism_overrides:atmosphere.delta_P.reference_year_doc = "Reference year to use when ``atmosphere.delta_P.period`` is active.";
    pism_overrides:atmosphere.delta_P.reference_year_option = "atmosphere_delta_P_reference_year";
    pism_overrides:atmosphere.delta_P.reference_year_type = "integer";
    pism_overrides:atmosphere.delta_P.reference_year_units = "years";

    pism_overrides:atmosphere.delta_T.file = "";
    pism_overrides:atmosphere.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_overrides:atmosphere.delta_T.file_option = "atmosphere_delta_T_file";
    pism_overrides:atmosphere.delta_T.file_type = "string";

    pism_overrides:atmosphere.delta_T.period = 0;
    pism_overrides:atmosphere.delta_T.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.delta_T.period_option = "atmosphere_delta_T_period";
    pism_overrides:atmosphere.delta_T.period_type = "integer";
    pism_overrides:atmosphere.delta_T.period_units = "years";

    pism_overrides:atmosphere.delta_T.reference_year = 0;
    pism_overrides:atmosphere.delta_T.reference_year_doc = "Reference year to use when ``atmosphere.delta_T.period`` is active.";
    pism_overrides:atmosphere.delta_T.reference_year_option = "atmosphere_delta_T_reference_year";
    pism_overrides:atmosphere.delta_T.reference_year_type = "integer";
    pism_overrides:atmosphere.delta_T.reference_year_units = "years";

    pism_overrides:atmosphere.elevation_change.file = "";
    pism_overrides:atmosphere.elevation_change.file_doc = "Name of the file containing the reference surface elevation field (variable ``usurf``).";
    pism_overrides:atmosphere.elevation_change.file_option = "atmosphere_lapse_rate_file";
    pism_overrides:atmosphere.elevation_change.file_type = "string";

    pism_overrides:atmosphere.elevation_change.period = 0;
    pism_overrides:atmosphere.elevation_change.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.elevation_change.period_option = "atmosphere_lapse_rate_period";
    pism_overrides:atmosphere.elevation_change.period_type = "integer";
    pism_overrides:atmosphere.elevation_change.period_units = "years";

    pism_overrides:atmosphere.elevation_change.precipitation.lapse_rate = 0.0;
    pism_overrides:atmosphere.elevation_change.precipitation.lapse_rate_doc = "Elevation lapse rate for the surface mass balance";
    pism_overrides:atmosphere.elevation_change.precipitation.lapse_rate_option = "precip_lapse_rate";
    pism_overrides:atmosphere.elevation_change.precipitation.lapse_rate_type = "number";
    pism_overrides:atmosphere.elevation_change.precipitation.lapse_rate_units = "(kg m-2 / year) / km";

    pism_overrides:atmosphere.elevation_change.precipitation.method = "shift";
    pism_overrides:atmosphere.elevation_change.precipitation.method_choices = "scale,shift";
    pism_overrides:atmosphere.elevation_change.precipitation.method_doc = "Choose the precipitation adjustment method. ``scale``: use temperature-change-dependent scaling factor. ``shift``: use the precipitation lapse rate.";
    pism_overrides:atmosphere.elevation_change.precipitation.method_option = "precip_adjustment";
    pism_overrides:atmosphere.elevation_change.precipitation.method_type = "keyword";

    pism_overrides:atmosphere.elevation_change.reference_year = 0;
    pism_overrides:atmosphere.elevation_change.reference_year_doc = "Reference year to use when ``atmosphere.elevation_change.period`` is active.";
    pism_overrides:atmosphere.elevation_change.reference_year_option = "atmosphere_lapse_rate_reference_year";
    pism_overrides:atmosphere.elevation_change.reference_year_type = "integer";
    pism_overrides:atmosphere.elevation_change.reference_year_units = "years";

    pism_overrides:atmosphere.elevation_change.temperature_lapse_rate = 0.0;
    pism_overrides:atmosphere.elevation_change.temperature_lapse_rate_doc = "Elevation lapse rate for the surface temperature";
    pism_overrides:atmosphere.elevation_change.temperature_lapse_rate_option = "temp_lapse_rate";
    pism_overrides:atmosphere.elevation_change.temperature_lapse_rate_type = "number";
    pism_overrides:atmosphere.elevation_change.temperature_lapse_rate_units = "Kelvin / km";

    pism_overrides:atmosphere.fausto_air_temp.c_ma = -0.7189;
    pism_overrides:atmosphere.fausto_air_temp.c_ma_doc = "latitude-dependence coefficient for formula (1) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.c_ma_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.c_ma_units = "Kelvin / degree_north";

    pism_overrides:atmosphere.fausto_air_temp.c_mj = -0.1585;
    pism_overrides:atmosphere.fausto_air_temp.c_mj_doc = "latitude-dependence coefficient for formula (2) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.c_mj_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.c_mj_units = "Kelvin / degree_north";

    pism_overrides:atmosphere.fausto_air_temp.d_ma = 314.98;
    pism_overrides:atmosphere.fausto_air_temp.d_ma_doc = "41.83+273.15; base temperature for formula (1) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.d_ma_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.d_ma_units = "Kelvin";

    pism_overrides:atmosphere.fausto_air_temp.d_mj = 287.85;
    pism_overrides:atmosphere.fausto_air_temp.d_mj_doc = "= 14.70+273.15; base temperature for formula (2) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.d_mj_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.d_mj_units = "Kelvin";

    pism_overrides:atmosphere.fausto_air_temp.gamma_ma = -0.006309;
    pism_overrides:atmosphere.fausto_air_temp.gamma_ma_doc = "= -6.309 / 1km; mean slope lapse rate for formula (1) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.gamma_ma_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.gamma_ma_units = "Kelvin / meter";

    pism_overrides:atmosphere.fausto_air_temp.gamma_mj = -0.005426;
    pism_overrides:atmosphere.fausto_air_temp.gamma_mj_doc = "= -5.426 / 1km; mean slope lapse rate for formula (2) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.gamma_mj_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.gamma_mj_units = "Kelvin / meter";

    pism_overrides:atmosphere.fausto_air_temp.kappa_ma = 0.0672;
    pism_overrides:atmosphere.fausto_air_temp.kappa_ma_doc = "longitude-dependence coefficient for formula (1) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.kappa_ma_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.kappa_ma_units = "Kelvin / degree_west";

    pism_overrides:atmosphere.fausto_air_temp.kappa_mj = 0.0518;
    pism_overrides:atmosphere.fausto_air_temp.kappa_mj_doc = "longitude-dependence coefficient for formula (2) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.kappa_mj_type = "number";
    pism_overrides:atmosphere.fausto_air_temp.kappa_mj_units = "Kelvin / degree_west";

    pism_overrides:atmosphere.fausto_air_temp.summer_peak_day = 196;
    pism_overrides:atmosphere.fausto_air_temp.summer_peak_day_doc = "day of year for July 15; used in corrected formula (4) in :cite:`Faustoetal2009`";
    pism_overrides:atmosphere.fausto_air_temp.summer_peak_day_type = "integer";
    pism_overrides:atmosphere.fausto_air_temp.summer_peak_day_units = "ordinal day number";

    pism_overrides:atmosphere.frac_P.file = "";
    pism_overrides:atmosphere.frac_P.file_doc = "Name of the file containing scalar precipitation scaling.";
    pism_overrides:atmosphere.frac_P.file_option = "atmosphere_frac_P_file";
    pism_overrides:atmosphere.frac_P.file_type = "string";

    pism_overrides:atmosphere.frac_P.period = 0;
    pism_overrides:atmosphere.frac_P.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.frac_P.period_option = "atmosphere_frac_P_period";
    pism_overrides:atmosphere.frac_P.period_type = "integer";
    pism_overrides:atmosphere.frac_P.period_units = "years";

    pism_overrides:atmosphere.frac_P.reference_year = 0;
    pism_overrides:atmosphere.frac_P.reference_year_doc = "Reference year to use when ``atmosphere.frac_P.period`` is active.";
    pism_overrides:atmosphere.frac_P.reference_year_option = "atmosphere_frac_P_reference_year";
    pism_overrides:atmosphere.frac_P.reference_year_type = "integer";
    pism_overrides:atmosphere.frac_P.reference_year_units = "years";

    pism_overrides:atmosphere.given.file = "";
    pism_overrides:atmosphere.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:atmosphere.given.file_option = "atmosphere_given_file";
    pism_overrides:atmosphere.given.file_type = "string";

    pism_overrides:atmosphere.given.period = 0;
    pism_overrides:atmosphere.given.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.given.period_option = "atmosphere_given_period";
    pism_overrides:atmosphere.given.period_type = "integer";
    pism_overrides:atmosphere.given.period_units = "years";

    pism_overrides:atmosphere.given.reference_year = 0;
    pism_overrides:atmosphere.given.reference_year_doc = "Reference year to use when ``atmosphere.given.period`` is active.";
    pism_overrides:atmosphere.given.reference_year_option = "atmosphere_given_reference_year";
    pism_overrides:atmosphere.given.reference_year_type = "integer";
    pism_overrides:atmosphere.given.reference_year_units = "years";

    pism_overrides:atmosphere.models = "given";
    pism_overrides:atmosphere.models_doc = "Comma-separated list of atmosphere melt models and modifiers.";
    pism_overrides:atmosphere.models_option = "atmosphere";
    pism_overrides:atmosphere.models_type = "string";

    pism_overrides:atmosphere.one_station.file = "";
    pism_overrides:atmosphere.one_station.file_doc = "Specifies a file containing scalar time-series 'precipitation' and 'air_temp'.";
    pism_overrides:atmosphere.one_station.file_option = "atmosphere_one_station_file";
    pism_overrides:atmosphere.one_station.file_type = "string";

    pism_overrides:atmosphere.orographic_precipitation.background_precip_post = 0;
    pism_overrides:atmosphere.orographic_precipitation.background_precip_post_doc = "Adding background precipitation after truncation";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_post_option = "background_precip_post";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_post_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_post_units = "mm/hr";

    pism_overrides:atmosphere.orographic_precipitation.background_precip_pre = 0;
    pism_overrides:atmosphere.orographic_precipitation.background_precip_pre_doc = "Adding background precipitation before truncation";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_pre_option = "background_precip_pre";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_pre_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.background_precip_pre_units = "mm/hr";

    pism_overrides:atmosphere.orographic_precipitation.conversion_time = 1000.0;
    pism_overrides:atmosphere.orographic_precipitation.conversion_time_doc = "Cloud conversion time";
    pism_overrides:atmosphere.orographic_precipitation.conversion_time_option = "conversion_time";
    pism_overrides:atmosphere.orographic_precipitation.conversion_time_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.conversion_time_units = "s";

    pism_overrides:atmosphere.orographic_precipitation.coriolis_latitude = 0.0;
    pism_overrides:atmosphere.orographic_precipitation.coriolis_latitude_doc = "Latitude used to compute Coriolis force";
    pism_overrides:atmosphere.orographic_precipitation.coriolis_latitude_option = "coriolis_latitude";
    pism_overrides:atmosphere.orographic_precipitation.coriolis_latitude_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.coriolis_latitude_units = "degrees_N";

    pism_overrides:atmosphere.orographic_precipitation.fallout_time = 1000.0;
    pism_overrides:atmosphere.orographic_precipitation.fallout_time_doc = "Fallout time";
    pism_overrides:atmosphere.orographic_precipitation.fallout_time_option = "fallout_time";
    pism_overrides:atmosphere.orographic_precipitation.fallout_time_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.fallout_time_units = "s";

    pism_overrides:atmosphere.orographic_precipitation.grid_size_factor = 2;
    pism_overrides:atmosphere.orographic_precipitation.grid_size_factor_doc = "The spectral grid size is (Z*(grid.Mx - 1) + 1, Z*(grid.My - 1) + 1) where Z is given by this parameter.";
    pism_overrides:atmosphere.orographic_precipitation.grid_size_factor_type = "integer";
    pism_overrides:atmosphere.orographic_precipitation.grid_size_factor_units = "count";

    pism_overrides:atmosphere.orographic_precipitation.lapse_rate = -5.8;
    pism_overrides:atmosphere.orographic_precipitation.lapse_rate_doc = "Lapse rate";
    pism_overrides:atmosphere.orographic_precipitation.lapse_rate_option = "lapse_rate";
    pism_overrides:atmosphere.orographic_precipitation.lapse_rate_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.lapse_rate_units = "K / km";

    pism_overrides:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate = -6.5;
    pism_overrides:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_doc = "Water vapor scale height";
    pism_overrides:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_option = "moist_adiabatic_lapse_rate";
    pism_overrides:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_units = "K / km";

    pism_overrides:atmosphere.orographic_precipitation.moist_stability_frequency = 0.05;
    pism_overrides:atmosphere.orographic_precipitation.moist_stability_frequency_doc = "Moist stability frequency";
    pism_overrides:atmosphere.orographic_precipitation.moist_stability_frequency_option = "moist_stability_frequency";
    pism_overrides:atmosphere.orographic_precipitation.moist_stability_frequency_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.moist_stability_frequency_units = "1/s";

    pism_overrides:atmosphere.orographic_precipitation.reference_density = 7.4e-3;
    pism_overrides:atmosphere.orographic_precipitation.reference_density_doc = "Water vapor scale height";
    pism_overrides:atmosphere.orographic_precipitation.reference_density_option = "reference_density";
    pism_overrides:atmosphere.orographic_precipitation.reference_density_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.reference_density_units = "kg m-3";

    pism_overrides:atmosphere.orographic_precipitation.scale_factor = 1;
    pism_overrides:atmosphere.orographic_precipitation.scale_factor_doc = "Precipitation scaling factor";
    pism_overrides:atmosphere.orographic_precipitation.scale_factor_option = "scale_factor";
    pism_overrides:atmosphere.orographic_precipitation.scale_factor_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.scale_factor_units = "1";

    pism_overrides:atmosphere.orographic_precipitation.truncate = "true";
    pism_overrides:atmosphere.orographic_precipitation.truncate_doc = "Truncate precipitation at 0";
    pism_overrides:atmosphere.orographic_precipitation.truncate_option = "truncate";
    pism_overrides:atmosphere.orographic_precipitation.truncate_type = "flag";

    pism_overrides:atmosphere.orographic_precipitation.water_vapor_scale_height = 2500.0;
    pism_overrides:atmosphere.orographic_precipitation.water_vapor_scale_height_doc = "Water vapor scale height";
    pism_overrides:atmosphere.orographic_precipitation.water_vapor_scale_height_option = "water_vapor_scale_height";
    pism_overrides:atmosphere.orographic_precipitation.water_vapor_scale_height_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.water_vapor_scale_height_units = "m";

    pism_overrides:atmosphere.orographic_precipitation.wind_direction = 270;
    pism_overrides:atmosphere.orographic_precipitation.wind_direction_doc = "The direction the wind is coming from";
    pism_overrides:atmosphere.orographic_precipitation.wind_direction_option = "wind_direction";
    pism_overrides:atmosphere.orographic_precipitation.wind_direction_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.wind_direction_units = "degrees";

    pism_overrides:atmosphere.orographic_precipitation.wind_speed = 10;
    pism_overrides:atmosphere.orographic_precipitation.wind_speed_doc = "The direction the wind is coming from";
    pism_overrides:atmosphere.orographic_precipitation.wind_speed_option = "wind_speed";
    pism_overrides:atmosphere.orographic_precipitation.wind_speed_type = "number";
    pism_overrides:atmosphere.orographic_precipitation.wind_speed_units = "m/s";

    pism_overrides:atmosphere.pik.file = "";
    pism_overrides:atmosphere.pik.file_doc = "Name of the file containing the reference surface elevation field (variable ``usurf``).";
    pism_overrides:atmosphere.pik.file_option = "atmosphere_pik_file";
    pism_overrides:atmosphere.pik.file_type = "string";

    pism_overrides:atmosphere.pik.parameterization = "martin";
    pism_overrides:atmosphere.pik.parameterization_choices = "martin,huybrechts_dewolde,martin_huybrechts_dewolde,era_interim,era_interim_sin,era_interim_lon";
    pism_overrides:atmosphere.pik.parameterization_doc = "Selects parameterizations of mean annual and mean summer near-surface air temperatures.";
    pism_overrides:atmosphere.pik.parameterization_option = "atmosphere_pik";
    pism_overrides:atmosphere.pik.parameterization_type = "keyword";

    pism_overrides:atmosphere.precip_exponential_factor_for_temperature = 0.07041666667;
    pism_overrides:atmosphere.precip_exponential_factor_for_temperature_doc = "= 0.169/2.4; in SeaRISE-Greenland formula for precipitation correction using air temperature offsets relative to present; a 7.3\% change of precipitation rate for every one degC of temperature change :cite:`Huybrechts02`";
    pism_overrides:atmosphere.precip_exponential_factor_for_temperature_type = "number";
    pism_overrides:atmosphere.precip_exponential_factor_for_temperature_units = "Kelvin-1";

    pism_overrides:atmosphere.precip_scaling.file = "";
    pism_overrides:atmosphere.precip_scaling.file_doc = "Name of the file containing temperature offsets to use for a precipitation correction.";
    pism_overrides:atmosphere.precip_scaling.file_option = "atmosphere_precip_scaling_file";
    pism_overrides:atmosphere.precip_scaling.file_type = "string";

    pism_overrides:atmosphere.precip_scaling.period = 0;
    pism_overrides:atmosphere.precip_scaling.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.precip_scaling.period_option = "atmosphere_precip_scaling_period";
    pism_overrides:atmosphere.precip_scaling.period_type = "integer";
    pism_overrides:atmosphere.precip_scaling.period_units = "years";

    pism_overrides:atmosphere.precip_scaling.reference_year = 0;
    pism_overrides:atmosphere.precip_scaling.reference_year_doc = "Reference year to use when ``atmosphere.precip_scaling.period`` is active.";
    pism_overrides:atmosphere.precip_scaling.reference_year_option = "atmosphere_precip_scaling_reference_year";
    pism_overrides:atmosphere.precip_scaling.reference_year_type = "integer";
    pism_overrides:atmosphere.precip_scaling.reference_year_units = "years";

    pism_overrides:atmosphere.searise_greenland.file = "";
    pism_overrides:atmosphere.searise_greenland.file_doc = "Name of the file containing a precipitation field.";
    pism_overrides:atmosphere.searise_greenland.file_option = "atmosphere_searise_greenland_file";
    pism_overrides:atmosphere.searise_greenland.file_type = "string";

    pism_overrides:atmosphere.uniform.precipitation = 1000;
    pism_overrides:atmosphere.uniform.precipitation_doc = "Precipitation used by the 'uniform' atmosphere model.";
    pism_overrides:atmosphere.uniform.precipitation_type = "number";
    pism_overrides:atmosphere.uniform.precipitation_units = "kg m-2 year-1";

    pism_overrides:atmosphere.uniform.temperature = 273.15;
    pism_overrides:atmosphere.uniform.temperature_doc = "Air temperature used by the 'uniform' atmosphere model.";
    pism_overrides:atmosphere.uniform.temperature_type = "number";
    pism_overrides:atmosphere.uniform.temperature_units = "Kelvin";

    pism_overrides:atmosphere.yearly_cycle.file = "";
    pism_overrides:atmosphere.yearly_cycle.file_doc = "Name of the file containing mean annual and mean July temperatures (`air_temp_mean_annual` and `air_temp_mean_summer`) and the `precipitation` field.";
    pism_overrides:atmosphere.yearly_cycle.file_option = "atmosphere_yearly_cycle_file";
    pism_overrides:atmosphere.yearly_cycle.file_type = "string";

    pism_overrides:atmosphere.yearly_cycle.scaling.file = "";
    pism_overrides:atmosphere.yearly_cycle.scaling.file_doc = "Name of the file containing amplitude scaling (`amplitude_scaling`) for the near-surface air temperature.";
    pism_overrides:atmosphere.yearly_cycle.scaling.file_option = "atmosphere_yearly_cycle_scaling_file";
    pism_overrides:atmosphere.yearly_cycle.scaling.file_type = "string";

    pism_overrides:atmosphere.yearly_cycle.scaling.period = 0;
    pism_overrides:atmosphere.yearly_cycle.scaling.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:atmosphere.yearly_cycle.scaling.period_type = "integer";
    pism_overrides:atmosphere.yearly_cycle.scaling.period_units = "years";

    pism_overrides:atmosphere.yearly_cycle.scaling.reference_year = 0;
    pism_overrides:atmosphere.yearly_cycle.scaling.reference_year_doc = "Reference year to use when ``atmosphere.yearly_cycle.scaling.period`` is active.";
    pism_overrides:atmosphere.yearly_cycle.scaling.reference_year_type = "integer";
    pism_overrides:atmosphere.yearly_cycle.scaling.reference_year_units = "years";

    pism_overrides:basal_resistance.beta_ice_free_bedrock = 1.8e9;
    pism_overrides:basal_resistance.beta_ice_free_bedrock_doc = "value is for ice stream E from :cite:`HulbeMacAyeal`; thus sliding velocity, but we hope it doesn't matter much; at 100 m/year the linear sliding law gives 57040 Pa basal shear stress";
    pism_overrides:basal_resistance.beta_ice_free_bedrock_type = "number";
    pism_overrides:basal_resistance.beta_ice_free_bedrock_units = "Pascal second meter-1";

    pism_overrides:basal_resistance.beta_lateral_margin = 1e19;
    pism_overrides:basal_resistance.beta_lateral_margin_doc = "high value of `\\beta` used to simulate drag at lateral ice margins (fjord walls, etc); the default value is chosen to disable flow in the direction along a margin";
    pism_overrides:basal_resistance.beta_lateral_margin_type = "number";
    pism_overrides:basal_resistance.beta_lateral_margin_units = "Pascal second meter-1";

    pism_overrides:basal_resistance.plastic.regularization = 0.01;
    pism_overrides:basal_resistance.plastic.regularization_doc = "Set the value of `\\epsilon` regularization of plastic till; this is the second `\\epsilon` in formula (4.1) in :cite:`SchoofStream`";
    pism_overrides:basal_resistance.plastic.regularization_option = "plastic_reg";
    pism_overrides:basal_resistance.plastic.regularization_type = "number";
    pism_overrides:basal_resistance.plastic.regularization_units = "meter / year";

    pism_overrides:basal_resistance.pseudo_plastic.enabled = "no";
    pism_overrides:basal_resistance.pseudo_plastic.enabled_doc = "Use the pseudo-plastic till model (basal sliding law).";
    pism_overrides:basal_resistance.pseudo_plastic.enabled_option = "pseudo_plastic";
    pism_overrides:basal_resistance.pseudo_plastic.enabled_type = "flag";

    pism_overrides:basal_resistance.pseudo_plastic.q = 0.25;
    pism_overrides:basal_resistance.pseudo_plastic.q_doc = "The exponent of the pseudo-plastic basal resistance model";
    pism_overrides:basal_resistance.pseudo_plastic.q_option = "pseudo_plastic_q";
    pism_overrides:basal_resistance.pseudo_plastic.q_type = "number";
    pism_overrides:basal_resistance.pseudo_plastic.q_units = "pure number";

    pism_overrides:basal_resistance.pseudo_plastic.sliding_scale_factor = -1.0;
    pism_overrides:basal_resistance.pseudo_plastic.sliding_scale_factor_doc = "divides pseudo-plastic tauc (yield stress) by given factor; this would increase sliding by given factor in absence of membrane stresses; not used if negative or zero; not used by default";
    pism_overrides:basal_resistance.pseudo_plastic.sliding_scale_factor_option = "sliding_scale_factor_reduces_tauc";
    pism_overrides:basal_resistance.pseudo_plastic.sliding_scale_factor_type = "number";
    pism_overrides:basal_resistance.pseudo_plastic.sliding_scale_factor_units = "1";

    pism_overrides:basal_resistance.pseudo_plastic.u_threshold = 100.0;
    pism_overrides:basal_resistance.pseudo_plastic.u_threshold_doc = "threshold velocity of the pseudo-plastic sliding law";
    pism_overrides:basal_resistance.pseudo_plastic.u_threshold_option = "pseudo_plastic_uthreshold";
    pism_overrides:basal_resistance.pseudo_plastic.u_threshold_type = "number";
    pism_overrides:basal_resistance.pseudo_plastic.u_threshold_units = "meter / year";

    pism_overrides:basal_yield_stress.add_transportable_water = "no";
    pism_overrides:basal_yield_stress.add_transportable_water_doc = "If 'yes' then the water amount in the transport system is added to tillwat in determining tauc (in the Mohr-Coulomb relation).  Normally only the water in the till is used.";
    pism_overrides:basal_yield_stress.add_transportable_water_option = "tauc_add_transportable_water";
    pism_overrides:basal_yield_stress.add_transportable_water_type = "flag";

    pism_overrides:basal_yield_stress.constant.value = 2e5;
    pism_overrides:basal_yield_stress.constant.value_doc = "fill value for yield stress for basal till (plastic or pseudo-plastic model); note `2 \\times 10^5` Pa = 2 bar is quite strong and little sliding should occur";
    pism_overrides:basal_yield_stress.constant.value_option = "tauc";
    pism_overrides:basal_yield_stress.constant.value_type = "number";
    pism_overrides:basal_yield_stress.constant.value_units = "Pascal";

    pism_overrides:basal_yield_stress.ice_free_bedrock = 1e6;
    pism_overrides:basal_yield_stress.ice_free_bedrock_doc = "the 'high' yield stress value used in grounded ice-free areas.";
    pism_overrides:basal_yield_stress.ice_free_bedrock_option = "high_tauc";
    pism_overrides:basal_yield_stress.ice_free_bedrock_type = "number";
    pism_overrides:basal_yield_stress.ice_free_bedrock_units = "Pascal";

    pism_overrides:basal_yield_stress.model = "mohr_coulomb";
    pism_overrides:basal_yield_stress.model_choices = "constant,mohr_coulomb";
    pism_overrides:basal_yield_stress.model_doc = "The basal yield stress model to use when sliding is active.";
    pism_overrides:basal_yield_stress.model_option = "yield_stress";
    pism_overrides:basal_yield_stress.model_type = "keyword";

    pism_overrides:basal_yield_stress.mohr_coulomb.delta.file = "";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.file_doc = "Name of the file containing space- and time-dependent variable `mohr_coulomb_delta` to use instead of `basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden`.";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.file_option = "mohr_coulomb_delta_file";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.file_type = "string";

    pism_overrides:basal_yield_stress.mohr_coulomb.delta.period = 0;
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.period_doc = "Length of the period. Set to zero to disable.";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.period_option = "mohr_coulomb_delta_period";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.period_type = "integer";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.period_units = "years";

    pism_overrides:basal_yield_stress.mohr_coulomb.delta.reference_year = 0;
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.reference_year_doc = "Reference year to use when ``basal_yield_stress.mohr_coulomb.delta.period`` is active.";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.reference_year_option = "mohr_coulomb_delta_reference_year";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.reference_year_type = "integer";
    pism_overrides:basal_yield_stress.mohr_coulomb.delta.reference_year_units = "years";

    pism_overrides:basal_yield_stress.mohr_coulomb.tauc_to_phi.file = "";
    pism_overrides:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_doc = "File containing the basal yield stress field that should be used to recover the till friction angle distribution.";
    pism_overrides:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_option = "tauc_to_phi";
    pism_overrides:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_type = "string";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_cohesion = 0.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_cohesion_doc = "cohesion of till; = c_0 in most references; note Schoof uses zero but Paterson pp 168--169 gives range 0--40 kPa; but Paterson notes that '... all the pairs c_0 and phi in the table would give a yield stress for Ice Stream B that exceeds the basal shear stress there...'";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_cohesion_option = "till_cohesion";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_cohesion_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_cohesion_units = "Pascal";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient = 0.12;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_doc = "coefficient of compressiblity of till; value from :cite:`Tulaczyketal2000`";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_option = "till_compressibility_coefficient";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_units = "pure number";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden = 0.02;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_doc = "`\\delta` in notes; `N_0 = \\delta P_o` where `P_o` is overburden pressure; `N_0` is reference (low) value of effective pressure (i.e. normal stress); `N_0` scales with overburden pressure unlike :cite:`Tulaczyketal2000`; default value from Greenland and Antarctic model runs";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_option = "till_effective_fraction_overburden";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_units = "pure number";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water = 0.1;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_doc = "If basal_yield_stress.add_transportable_water = yes then the water amount in the transport system is added to tillwat in determining tauc.  Normally only the water in the till is used.  This factor multiplies the logarithm in that formula.";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_option = "till_log_factor_transportable_water";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_units = "meters";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_phi_default = 30.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_phi_default_doc = "fill value for till friction angle";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_phi_default_option = "plastic_phi";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_phi_default_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_phi_default_units = "degrees";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure = 1000.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_doc = "reference effective pressure N_0; value from :cite:`Tulaczyketal2000`";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_units = "Pascal";

    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_void_ratio = 0.69;
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_doc = "void ratio at reference effective pressure N_0; value from :cite:`Tulaczyketal2000`";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_option = "till_reference_void_ratio";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_units = "pure number";

    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled = "no";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_doc = "If the option ``-topg_to_phi`` is set then this will be set to 'yes', and then MohrCoulombYieldStress will initialize the ``tillphi`` field using a piece-wise linear function of depth described by four parameters.";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_type = "flag";

    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max = 15.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_doc = "upper value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_units = "degrees";

    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min = 5.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_doc = "lower value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_units = "degrees";

    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max = 1000.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_doc = "the elevation at which the upper value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_units = "meters";

    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min = -1000.0;
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_doc = "the elevation at which the lower value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_type = "number";
    pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_units = "meters";

    pism_overrides:basal_yield_stress.slippery_grounding_lines = "no";
    pism_overrides:basal_yield_stress.slippery_grounding_lines_doc = "If yes, at icy grounded locations with bed elevations below sea level, within one cell of floating ice or ice-free ocean, make tauc as low as possible from the Mohr-Coulomb relation.  Specifically, at such locations replace the normally-computed tauc from the Mohr-Coulomb relation, which uses the effective pressure from the modeled amount of water in the till, by the minimum value of tauc from Mohr-Coulomb, i.e. by using the effective pressure corresponding to the maximum amount of till-stored water.  Does not alter the modeled or reported amount of till water, nor does this mechanism affect water conservation.";
    pism_overrides:basal_yield_stress.slippery_grounding_lines_option = "tauc_slippery_grounding_lines";
    pism_overrides:basal_yield_stress.slippery_grounding_lines_type = "flag";

    pism_overrides:bed_deformation.bed_topography_delta_file = "";
    pism_overrides:bed_deformation.bed_topography_delta_file_doc = "The name of the file to read the topg_delta from. This field is added to the bed topography during initialization.";
    pism_overrides:bed_deformation.bed_topography_delta_file_option = "topg_delta_file";
    pism_overrides:bed_deformation.bed_topography_delta_file_type = "string";

    pism_overrides:bed_deformation.bed_uplift_file = "";
    pism_overrides:bed_deformation.bed_uplift_file_doc = "The name of the file to read the uplift (dbdt) from. Leave empty to read it from an input file or a regridding file.";
    pism_overrides:bed_deformation.bed_uplift_file_option = "uplift_file";
    pism_overrides:bed_deformation.bed_uplift_file_type = "string";

    pism_overrides:bed_deformation.lc.elastic_model = "yes";
    pism_overrides:bed_deformation.lc.elastic_model_doc = "Use the elastic part of the Lingle-Clark bed deformation model.";
    pism_overrides:bed_deformation.lc.elastic_model_option = "bed_def_lc_elastic_model";
    pism_overrides:bed_deformation.lc.elastic_model_type = "flag";

    pism_overrides:bed_deformation.lc.grid_size_factor = 4;
    pism_overrides:bed_deformation.lc.grid_size_factor_doc = "The spectral grid size is (Z*(grid.Mx - 1) + 1, Z*(grid.My - 1) + 1) where Z is given by this parameter. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_overrides:bed_deformation.lc.grid_size_factor_type = "integer";
    pism_overrides:bed_deformation.lc.grid_size_factor_units = "count";

    pism_overrides:bed_deformation.lc.update_interval = 10.0;
    pism_overrides:bed_deformation.lc.update_interval_doc = "Interval between updates of the Lingle-Clark model";
    pism_overrides:bed_deformation.lc.update_interval_type = "number";
    pism_overrides:bed_deformation.lc.update_interval_units = "years";

    pism_overrides:bed_deformation.lithosphere_flexural_rigidity = 5.0e24;
    pism_overrides:bed_deformation.lithosphere_flexural_rigidity_doc = "lithosphere flexural rigidity used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_overrides:bed_deformation.lithosphere_flexural_rigidity_type = "number";
    pism_overrides:bed_deformation.lithosphere_flexural_rigidity_units = "Newton meter";

    pism_overrides:bed_deformation.mantle_density = 3300.0;
    pism_overrides:bed_deformation.mantle_density_doc = "half-space (mantle) density used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_overrides:bed_deformation.mantle_density_type = "number";
    pism_overrides:bed_deformation.mantle_density_units = "kg meter-3";

    pism_overrides:bed_deformation.mantle_viscosity = 1.0e21;
    pism_overrides:bed_deformation.mantle_viscosity_doc = "half-space (mantle) viscosity used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_overrides:bed_deformation.mantle_viscosity_type = "number";
    pism_overrides:bed_deformation.mantle_viscosity_units = "Pascal second";

    pism_overrides:bed_deformation.model = "none";
    pism_overrides:bed_deformation.model_choices = "none,iso,lc";
    pism_overrides:bed_deformation.model_doc = "Selects a bed deformation model to use. 'iso' is point-wise isostasy, 'lc' is the Lingle-Clark model (see :cite:`LingleClark`, requires FFTW3).";
    pism_overrides:bed_deformation.model_option = "bed_def";
    pism_overrides:bed_deformation.model_type = "keyword";

    pism_overrides:bootstrapping.defaults.bed = 1.0;
    pism_overrides:bootstrapping.defaults.bed_doc = "bed elevation value to use if topg (bedrock_altitude) variable is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.bed_type = "number";
    pism_overrides:bootstrapping.defaults.bed_units = "meters";

    pism_overrides:bootstrapping.defaults.bmelt = 0.0;
    pism_overrides:bootstrapping.defaults.bmelt_doc = "basal melt rate value to use if variable bmelt is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.bmelt_type = "number";
    pism_overrides:bootstrapping.defaults.bmelt_units = "meter / second";

    pism_overrides:bootstrapping.defaults.bwat = 0.0;
    pism_overrides:bootstrapping.defaults.bwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.bwat_type = "number";
    pism_overrides:bootstrapping.defaults.bwat_units = "meters";

    pism_overrides:bootstrapping.defaults.bwp = 0.0;
    pism_overrides:bootstrapping.defaults.bwp_doc = "basal water pressure value to use if variable bwp is absent in bootstrapping file; most hydrology models do not use this value because bwp is diagnostic";
    pism_overrides:bootstrapping.defaults.bwp_type = "number";
    pism_overrides:bootstrapping.defaults.bwp_units = "Pascal";

    pism_overrides:bootstrapping.defaults.enwat = 0.0;
    pism_overrides:bootstrapping.defaults.enwat_doc = "effective englacial water thickness value to use if variable enwat is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.enwat_type = "number";
    pism_overrides:bootstrapping.defaults.enwat_units = "meters";

    pism_overrides:bootstrapping.defaults.geothermal_flux = 0.042;
    pism_overrides:bootstrapping.defaults.geothermal_flux_doc = "geothermal flux value to use if bheatflx variable is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.geothermal_flux_type = "number";
    pism_overrides:bootstrapping.defaults.geothermal_flux_units = "Watt meter-2";

    pism_overrides:bootstrapping.defaults.ice_thickness = 0.0;
    pism_overrides:bootstrapping.defaults.ice_thickness_doc = "thickness value to use if thk (land_ice_thickness) variable is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.ice_thickness_type = "number";
    pism_overrides:bootstrapping.defaults.ice_thickness_units = "meters";

    pism_overrides:bootstrapping.defaults.tillwat = 0.0;
    pism_overrides:bootstrapping.defaults.tillwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.tillwat_type = "number";
    pism_overrides:bootstrapping.defaults.tillwat_units = "meters";

    pism_overrides:bootstrapping.defaults.uplift = 0.0;
    pism_overrides:bootstrapping.defaults.uplift_doc = "uplift value to use if dbdt variable is absent in bootstrapping file";
    pism_overrides:bootstrapping.defaults.uplift_type = "number";
    pism_overrides:bootstrapping.defaults.uplift_units = "meter / second";

    pism_overrides:bootstrapping.temperature_heuristic = "smb";
    pism_overrides:bootstrapping.temperature_heuristic_choices = "smb,quartic_guess";
    pism_overrides:bootstrapping.temperature_heuristic_doc = "The heuristic to use to initialize ice temperature during bootstrapping: 'smb' uses the surface mass balance, surface temperature, and the geothermal flux, 'quartic_guess' uses the surface temperature and the geothermal flux.";
    pism_overrides:bootstrapping.temperature_heuristic_option = "boot_temperature_heuristic";
    pism_overrides:bootstrapping.temperature_heuristic_type = "keyword";

    pism_overrides:calving.eigen_calving.K = 0.0;
    pism_overrides:calving.eigen_calving.K_doc = "Set proportionality constant to determine calving rate from strain rates.  Note references :cite:`Levermannetal2012`, :cite:`Martinetal2011` use K in range `10^{9}` to `3 \\times 10^{11}` m a, that is, `3 \\times 10^{16}` to `10^{19}` m s.";
    pism_overrides:calving.eigen_calving.K_option = "eigen_calving_K";
    pism_overrides:calving.eigen_calving.K_type = "number";
    pism_overrides:calving.eigen_calving.K_units = "meter second";

    pism_overrides:calving.float_kill.calve_near_grounding_line = "yes";
    pism_overrides:calving.float_kill.calve_near_grounding_line_doc = "Calve floating ice near the grounding line.";
    pism_overrides:calving.float_kill.calve_near_grounding_line_option = "float_kill_calve_near_grounding_line";
    pism_overrides:calving.float_kill.calve_near_grounding_line_type = "flag";

    pism_overrides:calving.float_kill.margin_only = "no";
    pism_overrides:calving.float_kill.margin_only_doc = "Apply float_kill at ice margin cells only.";
    pism_overrides:calving.float_kill.margin_only_option = "float_kill_margin_only";
    pism_overrides:calving.float_kill.margin_only_type = "flag";

    pism_overrides:calving.hayhurst_calving.B_tilde = 65.0;
    pism_overrides:calving.hayhurst_calving.B_tilde_doc = "Effective damage rate :cite:`Mercenier2018`";
    pism_overrides:calving.hayhurst_calving.B_tilde_type = "number";
    pism_overrides:calving.hayhurst_calving.B_tilde_units = "(MPa)^r / year";

    pism_overrides:calving.hayhurst_calving.exponent_r = 0.43;
    pism_overrides:calving.hayhurst_calving.exponent_r_doc = "Damage law exponent :cite:`Mercenier2018`";
    pism_overrides:calving.hayhurst_calving.exponent_r_type = "number";
    pism_overrides:calving.hayhurst_calving.exponent_r_units = "1";

    pism_overrides:calving.hayhurst_calving.sigma_threshold = 0.17;
    pism_overrides:calving.hayhurst_calving.sigma_threshold_doc = "Damage threshold stress :cite:`Mercenier2018`";
    pism_overrides:calving.hayhurst_calving.sigma_threshold_type = "number";
    pism_overrides:calving.hayhurst_calving.sigma_threshold_units = "MPa";

    pism_overrides:calving.methods = "";
    pism_overrides:calving.methods_doc = "comma-separated list of calving methods; one or more of 'eigen_calving', 'float_kill', 'thickness_calving'";
    pism_overrides:calving.methods_option = "calving";
    pism_overrides:calving.methods_type = "string";

    pism_overrides:calving.thickness_calving.threshold = 50.0;
    pism_overrides:calving.thickness_calving.threshold_doc = "When terminal ice thickness of floating ice shelf is less than this threshold, it will be calved off.";
    pism_overrides:calving.thickness_calving.threshold_option = "thickness_calving_threshold";
    pism_overrides:calving.thickness_calving.threshold_type = "number";
    pism_overrides:calving.thickness_calving.threshold_units = "meters";

    pism_overrides:calving.thickness_calving.threshold_file = "";
    pism_overrides:calving.thickness_calving.threshold_file_doc = "Name of the file containing the spatially-variable thickness calving threshold.";
    pism_overrides:calving.thickness_calving.threshold_file_option = "thickness_calving_threshold_file";
    pism_overrides:calving.thickness_calving.threshold_file_type = "string";

    pism_overrides:calving.vonmises_calving.Glen_exponent = 3.0;
    pism_overrides:calving.vonmises_calving.Glen_exponent_doc = "Glen exponent in ice flow law for von Mises calving";
    pism_overrides:calving.vonmises_calving.Glen_exponent_option = "vonmises_calving_n";
    pism_overrides:calving.vonmises_calving.Glen_exponent_type = "number";
    pism_overrides:calving.vonmises_calving.Glen_exponent_units = "pure number";

    pism_overrides:calving.vonmises_calving.enhancement_factor = 1.0;
    pism_overrides:calving.vonmises_calving.enhancement_factor_doc = "Flow enhancement factor used by the flow law in the von Mises stress computation";
    pism_overrides:calving.vonmises_calving.enhancement_factor_type = "number";
    pism_overrides:calving.vonmises_calving.enhancement_factor_units = "1";

    pism_overrides:calving.vonmises_calving.enhancement_factor_interglacial = 1.0;
    pism_overrides:calving.vonmises_calving.enhancement_factor_interglacial_doc = "Flow enhancement factor used by the flow law in the von Mises stress computation (for ice accumulated during interglacial periods).";
    pism_overrides:calving.vonmises_calving.enhancement_factor_interglacial_type = "number";
    pism_overrides:calving.vonmises_calving.enhancement_factor_interglacial_units = "1";

    pism_overrides:calving.vonmises_calving.flow_law = "gpbld";
    pism_overrides:calving.vonmises_calving.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb";
    pism_overrides:calving.vonmises_calving.flow_law_doc = "The custom flow law for the von Mises stress computation";
    pism_overrides:calving.vonmises_calving.flow_law_type = "keyword";

    pism_overrides:calving.vonmises_calving.sigma_max = 1.0e6;
    pism_overrides:calving.vonmises_calving.sigma_max_doc = "Set maximum tensile stress.  Note references :cite:`Morlighem2016` use 1.0e6 Pa.";
    pism_overrides:calving.vonmises_calving.sigma_max_option = "vonmises_calving_calving_sigma_max";
    pism_overrides:calving.vonmises_calving.sigma_max_type = "number";
    pism_overrides:calving.vonmises_calving.sigma_max_units = "Pa";

    pism_overrides:calving.vonmises_calving.threshold_file = "";
    pism_overrides:calving.vonmises_calving.threshold_file_doc = "Name of the file containing the spatially-variable vonmises_calving calving threshold.";
    pism_overrides:calving.vonmises_calving.threshold_file_option = "vonmises_calving_threshold_file";
    pism_overrides:calving.vonmises_calving.threshold_file_type = "string";

    pism_overrides:calving.vonmises_calving.use_custom_flow_law = "no";
    pism_overrides:calving.vonmises_calving.use_custom_flow_law_doc = "Use custom flow law in the von Mises stress computation";
    pism_overrides:calving.vonmises_calving.use_custom_flow_law_option = "vonmises_calving_use_custom_flow_law";
    pism_overrides:calving.vonmises_calving.use_custom_flow_law_type = "flag";

    pism_overrides:constants.fresh_water.density = 1000.0;
    pism_overrides:constants.fresh_water.density_doc = "density of fresh water";
    pism_overrides:constants.fresh_water.density_type = "number";
    pism_overrides:constants.fresh_water.density_units = "kg meter-3";

    pism_overrides:constants.fresh_water.latent_heat_of_fusion = 3.34e5;
    pism_overrides:constants.fresh_water.latent_heat_of_fusion_doc = "latent heat of fusion for water :cite:`AschwandenBlatter`";
    pism_overrides:constants.fresh_water.latent_heat_of_fusion_type = "number";
    pism_overrides:constants.fresh_water.latent_heat_of_fusion_units = "Joule / kg";

    pism_overrides:constants.fresh_water.melting_point_temperature = 273.15;
    pism_overrides:constants.fresh_water.melting_point_temperature_doc = "melting point of pure water";
    pism_overrides:constants.fresh_water.melting_point_temperature_type = "number";
    pism_overrides:constants.fresh_water.melting_point_temperature_units = "Kelvin";

    pism_overrides:constants.fresh_water.specific_heat_capacity = 4170.0;
    pism_overrides:constants.fresh_water.specific_heat_capacity_doc = "at melting point T_0 :cite:`AschwandenBlatter`";
    pism_overrides:constants.fresh_water.specific_heat_capacity_type = "number";
    pism_overrides:constants.fresh_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_overrides:constants.global_ocean_area = 3.625e14;
    pism_overrides:constants.global_ocean_area_doc = "area of the global ocean :cite:`Cogley2011`";
    pism_overrides:constants.global_ocean_area_type = "number";
    pism_overrides:constants.global_ocean_area_units = "meter2";

    pism_overrides:constants.ice.beta_Clausius_Clapeyron = 7.9e-8;
    pism_overrides:constants.ice.beta_Clausius_Clapeyron_doc = "Clausius-Clapeyron constant relating melting temperature and pressure: `\\beta = dT / dP` :cite:`Luethi2002`";
    pism_overrides:constants.ice.beta_Clausius_Clapeyron_type = "number";
    pism_overrides:constants.ice.beta_Clausius_Clapeyron_units = "Kelvin / Pascal";

    pism_overrides:constants.ice.density = 910.0;
    pism_overrides:constants.ice.density_doc = "`\\rho_i`; density of ice in ice sheet";
    pism_overrides:constants.ice.density_type = "number";
    pism_overrides:constants.ice.density_units = "kg meter-3";

    pism_overrides:constants.ice.grain_size = 1.0;
    pism_overrides:constants.ice.grain_size_doc = "Default constant ice grain size to use with the Goldsby-Kohlstedt :cite:`GoldsbyKohlstedt` flow law";
    pism_overrides:constants.ice.grain_size_option = "ice_grain_size";
    pism_overrides:constants.ice.grain_size_type = "number";
    pism_overrides:constants.ice.grain_size_units = "mm";

    pism_overrides:constants.ice.specific_heat_capacity = 2009.0;
    pism_overrides:constants.ice.specific_heat_capacity_doc = "specific heat capacity of pure ice at melting point T_0";
    pism_overrides:constants.ice.specific_heat_capacity_type = "number";
    pism_overrides:constants.ice.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_overrides:constants.ice.thermal_conductivity = 2.10;
    pism_overrides:constants.ice.thermal_conductivity_doc = "= W m-1 K-1; thermal conductivity of pure ice";
    pism_overrides:constants.ice.thermal_conductivity_type = "number";
    pism_overrides:constants.ice.thermal_conductivity_units = "Joule / (meter Kelvin second)";

    pism_overrides:constants.ideal_gas_constant = 8.31441;
    pism_overrides:constants.ideal_gas_constant_doc = "ideal gas constant";
    pism_overrides:constants.ideal_gas_constant_type = "number";
    pism_overrides:constants.ideal_gas_constant_units = "Joule / (mol Kelvin)";

    pism_overrides:constants.sea_water.density = 1028.0;
    pism_overrides:constants.sea_water.density_doc = "density of sea water";
    pism_overrides:constants.sea_water.density_type = "number";
    pism_overrides:constants.sea_water.density_units = "kg meter-3";

    pism_overrides:constants.sea_water.specific_heat_capacity = 3985.0;
    pism_overrides:constants.sea_water.specific_heat_capacity_doc = "at 35 psu, value taken from `Kaye and Laby`_, section 2.7.9";
    pism_overrides:constants.sea_water.specific_heat_capacity_type = "number";
    pism_overrides:constants.sea_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_overrides:constants.standard_gravity = 9.81;
    pism_overrides:constants.standard_gravity_doc = "acceleration due to gravity on Earth geoid";
    pism_overrides:constants.standard_gravity_type = "number";
    pism_overrides:constants.standard_gravity_units = "meter second-2";

    pism_overrides:energy.allow_temperature_above_melting = "no";
    pism_overrides:energy.allow_temperature_above_melting_doc = "If set to 'yes', allow temperatures above the pressure-malting point in the cold mode temperature code. Used by some verifiaction tests.";
    pism_overrides:energy.allow_temperature_above_melting_type = "flag";

    pism_overrides:energy.basal_melt.use_grounded_cell_fraction  = "true";
    pism_overrides:energy.basal_melt.use_grounded_cell_fraction_doc = "If geometry.grounded_cell_fraction is set, use the fractional floatation mask to interpolate the basal melt rate at the grounding line between grounded and floating values.";
    pism_overrides:energy.basal_melt.use_grounded_cell_fraction_option  = "subgl_basal_melt";
    pism_overrides:energy.basal_melt.use_grounded_cell_fraction_type  = "flag";

    pism_overrides:energy.bedrock_thermal.conductivity = 3.0;
    pism_overrides:energy.bedrock_thermal.conductivity_doc = "= W m-1 K-1; for bedrock used in thermal model :cite:`RitzEISMINT`";
    pism_overrides:energy.bedrock_thermal.conductivity_type = "number";
    pism_overrides:energy.bedrock_thermal.conductivity_units = "Joule / (meter Kelvin second)";

    pism_overrides:energy.bedrock_thermal.density = 3300.0;
    pism_overrides:energy.bedrock_thermal.density_doc = "for bedrock used in thermal model";
    pism_overrides:energy.bedrock_thermal.density_type = "number";
    pism_overrides:energy.bedrock_thermal.density_units = "kg meter-3";

    pism_overrides:energy.bedrock_thermal.file = "";
    pism_overrides:energy.bedrock_thermal.file_doc = "Name of the file containing the geothermal flux field :var:`bheatflx`. Leave empty to read it from the :config:`input.file`.";
    pism_overrides:energy.bedrock_thermal.file_type = "string";

    pism_overrides:energy.bedrock_thermal.specific_heat_capacity = 1000.0;
    pism_overrides:energy.bedrock_thermal.specific_heat_capacity_doc = "for bedrock used in thermal model :cite:`RitzEISMINT`";
    pism_overrides:energy.bedrock_thermal.specific_heat_capacity_type = "number";
    pism_overrides:energy.bedrock_thermal.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_overrides:energy.ch_warming.average_channel_spacing = 20.0;
    pism_overrides:energy.ch_warming.average_channel_spacing_doc = "Average spacing between elements of the cryo-hydrologic system (controls the rate of heat transfer from the CH system into the ice).";
    pism_overrides:energy.ch_warming.average_channel_spacing_type = "number";
    pism_overrides:energy.ch_warming.average_channel_spacing_units = "meters";

    pism_overrides:energy.ch_warming.enabled = "no";
    pism_overrides:energy.ch_warming.enabled_doc = "Enable the cryo-hydrologic warming model";
    pism_overrides:energy.ch_warming.enabled_type = "flag";

    pism_overrides:energy.ch_warming.residual_water_fraction = 0.005;
    pism_overrides:energy.ch_warming.residual_water_fraction_doc = "residual water fraction in the cryo-hydrologic system at the end of a melt season";
    pism_overrides:energy.ch_warming.residual_water_fraction_type = "number";
    pism_overrides:energy.ch_warming.residual_water_fraction_units = "pure number";

    pism_overrides:energy.ch_warming.temperate_ice_thermal_conductivity_ratio = 1.0;
    pism_overrides:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_doc = "ratio of thermal conductivities of temperate and cold ice in the cryo-hydrologic system";
    pism_overrides:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_type = "number";
    pism_overrides:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_units = "pure number";

    pism_overrides:energy.drainage_maximum_rate = 1.58443823077064e-09;
    pism_overrides:energy.drainage_maximum_rate_doc = "0.05 year-1; maximum rate at which liquid water fraction in temperate ice could possibly drain; see :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_overrides:energy.drainage_maximum_rate_type = "number";
    pism_overrides:energy.drainage_maximum_rate_units = "second-1";

    pism_overrides:energy.drainage_target_water_fraction = 0.01;
    pism_overrides:energy.drainage_target_water_fraction_doc = "liquid water fraction (omega) above which drainage occurs, but below which there is no drainage; see :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_overrides:energy.drainage_target_water_fraction_type = "number";
    pism_overrides:energy.drainage_target_water_fraction_units = "1";

    pism_overrides:energy.enabled = "yes";
    pism_overrides:energy.enabled_doc = "Solve energy conservation equations.";
    pism_overrides:energy.enabled_type = "flag";

    pism_overrides:energy.enthalpy.cold_bulge_max = 60270.0;
    pism_overrides:energy.enthalpy.cold_bulge_max_doc = "= (2009 J kg-1 K-1) * (30 K); maximum amount by which advection can reduce the enthalpy of a column of ice below its surface enthalpy value";
    pism_overrides:energy.enthalpy.cold_bulge_max_type = "number";
    pism_overrides:energy.enthalpy.cold_bulge_max_units = "Joule / kg";

    pism_overrides:energy.enthalpy.temperate_ice_thermal_conductivity_ratio = 0.1;
    pism_overrides:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_doc = "K in cold ice is multiplied by this fraction to give K0 in :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_overrides:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_type = "number";
    pism_overrides:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_units = "pure number";

    pism_overrides:energy.margin_exclude_horizontal_advection = "yes";
    pism_overrides:energy.margin_exclude_horizontal_advection_doc = "Exclude horizontal advection of energy at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_overrides:energy.margin_exclude_horizontal_advection_type = "flag";

    pism_overrides:energy.margin_exclude_strain_heating = "yes";
    pism_overrides:energy.margin_exclude_strain_heating_doc = "Exclude strain heating at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_overrides:energy.margin_exclude_strain_heating_type = "flag";

    pism_overrides:energy.margin_exclude_vertical_advection = "yes";
    pism_overrides:energy.margin_exclude_vertical_advection_doc = "Exclude vertical advection of energy at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_overrides:energy.margin_exclude_vertical_advection_type = "flag";

    pism_overrides:energy.margin_ice_thickness_limit = 100.0;
    pism_overrides:energy.margin_ice_thickness_limit_doc = "use special margin treatment at grid points with a neighbor with the thickness below this limit.";
    pism_overrides:energy.margin_ice_thickness_limit_type = "number";
    pism_overrides:energy.margin_ice_thickness_limit_units = "meters";

    pism_overrides:energy.max_low_temperature_count = 10;
    pism_overrides:energy.max_low_temperature_count_doc = "Maximum number of grid points with ice temperature below energy.minimum_allowed_temperature.";
    pism_overrides:energy.max_low_temperature_count_option = "max_low_temps";
    pism_overrides:energy.max_low_temperature_count_type = "integer";
    pism_overrides:energy.max_low_temperature_count_units = "count";

    pism_overrides:energy.minimum_allowed_temperature = 200.0;
    pism_overrides:energy.minimum_allowed_temperature_doc = "Minimum allowed ice temperature";
    pism_overrides:energy.minimum_allowed_temperature_option = "low_temp";
    pism_overrides:energy.minimum_allowed_temperature_type = "number";
    pism_overrides:energy.minimum_allowed_temperature_units = "Kelvin";

    pism_overrides:energy.temperature_based = "no";
    pism_overrides:energy.temperature_based_doc = "Use cold ice (i.e. not polythermal) methods.";
    pism_overrides:energy.temperature_based_type = "flag";

    pism_overrides:energy.temperature_dependent_thermal_conductivity = "no";
    pism_overrides:energy.temperature_dependent_thermal_conductivity_doc = "If yes, use varkenthSystemCtx class in the energy step. It is base on formula (4.37) in :cite:`GreveBlatter2009`. Otherwise use enthSystemCtx, which has temperature-independent thermal conductivity set by constant ice.thermal_conductivity.";
    pism_overrides:energy.temperature_dependent_thermal_conductivity_option = "vark";
    pism_overrides:energy.temperature_dependent_thermal_conductivity_type = "flag";

    pism_overrides:enthalpy_converter.T_reference = 223.15;
    pism_overrides:enthalpy_converter.T_reference_doc = "= T_0 in enthalpy formulas in :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_overrides:enthalpy_converter.T_reference_type = "number";
    pism_overrides:enthalpy_converter.T_reference_units = "Kelvin";

    pism_overrides:enthalpy_converter.relaxed_is_temperate_tolerance = 0.001;
    pism_overrides:enthalpy_converter.relaxed_is_temperate_tolerance_doc = "Tolerance within which ice is treated as temperate (cold-ice mode and diagnostics).";
    pism_overrides:enthalpy_converter.relaxed_is_temperate_tolerance_type = "number";
    pism_overrides:enthalpy_converter.relaxed_is_temperate_tolerance_units = "Kelvin";

    pism_overrides:flow_law.Hooke.A = 4.42165e-9;
    pism_overrides:flow_law.Hooke.A_doc = "`A_{\\text{Hooke}} = (1/B_0)^n` where n=3 and B_0 = 1.928 `a^{1/3}` Pa. See :cite:`Hooke`";
    pism_overrides:flow_law.Hooke.A_type = "number";
    pism_overrides:flow_law.Hooke.A_units = "Pascal-3 second-1";

    pism_overrides:flow_law.Hooke.C = 0.16612;
    pism_overrides:flow_law.Hooke.C_doc = "See :cite:`Hooke`";
    pism_overrides:flow_law.Hooke.C_type = "number";
    pism_overrides:flow_law.Hooke.C_units = "Kelvin^{flow_law.Hooke.k}";

    pism_overrides:flow_law.Hooke.Q = 7.88e4;
    pism_overrides:flow_law.Hooke.Q_doc = "Activation energy, see :cite:`Hooke`";
    pism_overrides:flow_law.Hooke.Q_type = "number";
    pism_overrides:flow_law.Hooke.Q_units = "Joule / mol";

    pism_overrides:flow_law.Hooke.Tr = 273.39;
    pism_overrides:flow_law.Hooke.Tr_doc = "See :cite:`Hooke`";
    pism_overrides:flow_law.Hooke.Tr_type = "number";
    pism_overrides:flow_law.Hooke.Tr_units = "Kelvin";

    pism_overrides:flow_law.Hooke.k = 1.17;
    pism_overrides:flow_law.Hooke.k_doc = "See :cite:`Hooke`";
    pism_overrides:flow_law.Hooke.k_type = "number";
    pism_overrides:flow_law.Hooke.k_units = "pure number";

    pism_overrides:flow_law.Paterson_Budd.A_cold = 3.61e-13;
    pism_overrides:flow_law.Paterson_Budd.A_cold_doc = "Paterson-Budd A_cold, see :cite:`PatersonBudd`";
    pism_overrides:flow_law.Paterson_Budd.A_cold_type = "number";
    pism_overrides:flow_law.Paterson_Budd.A_cold_units = "Pascal-3 / second";

    pism_overrides:flow_law.Paterson_Budd.A_warm = 1.73e3;
    pism_overrides:flow_law.Paterson_Budd.A_warm_doc = "Paterson-Budd A_warm, see :cite:`PatersonBudd`";
    pism_overrides:flow_law.Paterson_Budd.A_warm_type = "number";
    pism_overrides:flow_law.Paterson_Budd.A_warm_units = "Pascal-3 / second";

    pism_overrides:flow_law.Paterson_Budd.Q_cold = 6.0e4;
    pism_overrides:flow_law.Paterson_Budd.Q_cold_doc = "Paterson-Budd Q_cold, see :cite:`PatersonBudd`";
    pism_overrides:flow_law.Paterson_Budd.Q_cold_type = "number";
    pism_overrides:flow_law.Paterson_Budd.Q_cold_units = "Joule / mol";

    pism_overrides:flow_law.Paterson_Budd.Q_warm = 13.9e4;
    pism_overrides:flow_law.Paterson_Budd.Q_warm_doc = "Paterson-Budd Q_warm, see :cite:`PatersonBudd`";
    pism_overrides:flow_law.Paterson_Budd.Q_warm_type = "number";
    pism_overrides:flow_law.Paterson_Budd.Q_warm_units = "Joule / mol";

    pism_overrides:flow_law.Paterson_Budd.T_critical = 263.15;
    pism_overrides:flow_law.Paterson_Budd.T_critical_doc = "Paterson-Budd critical temperature, see :cite:`PatersonBudd`";
    pism_overrides:flow_law.Paterson_Budd.T_critical_type = "number";
    pism_overrides:flow_law.Paterson_Budd.T_critical_units = "Kelvin";

    pism_overrides:flow_law.Schoof_regularizing_length = 1000.0;
    pism_overrides:flow_law.Schoof_regularizing_length_doc = "Regularizing length (Schoof definition)";
    pism_overrides:flow_law.Schoof_regularizing_length_type = "number";
    pism_overrides:flow_law.Schoof_regularizing_length_units = "km";

    pism_overrides:flow_law.Schoof_regularizing_velocity = 1.0;
    pism_overrides:flow_law.Schoof_regularizing_velocity_doc = "Regularizing velocity (Schoof definition)";
    pism_overrides:flow_law.Schoof_regularizing_velocity_type = "number";
    pism_overrides:flow_law.Schoof_regularizing_velocity_units = "meter / year";

    pism_overrides:flow_law.gpbld.water_frac_coeff = 181.25;
    pism_overrides:flow_law.gpbld.water_frac_coeff_doc = "coefficient in Glen-Paterson-Budd flow law for extra dependence of softness on liquid water fraction (omega) :cite:`GreveBlatter2009`, :cite:`LliboutryDuval1985`";
    pism_overrides:flow_law.gpbld.water_frac_coeff_type = "number";
    pism_overrides:flow_law.gpbld.water_frac_coeff_units = "pure number";

    pism_overrides:flow_law.gpbld.water_frac_observed_limit = 0.01;
    pism_overrides:flow_law.gpbld.water_frac_observed_limit_doc = "maximum value of liquid water fraction omega for which softness values are parameterized by :cite:`LliboutryDuval1985`; used in Glen-Paterson-Budd-Lliboutry-Duval flow law; compare :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_overrides:flow_law.gpbld.water_frac_observed_limit_type = "number";
    pism_overrides:flow_law.gpbld.water_frac_observed_limit_units = "1";

    pism_overrides:flow_law.isothermal_Glen.ice_softness = 3.1689e-24;
    pism_overrides:flow_law.isothermal_Glen.ice_softness_doc = "ice softness used by IsothermalGlenIce :cite:`EISMINT96`";
    pism_overrides:flow_law.isothermal_Glen.ice_softness_type = "number";
    pism_overrides:flow_law.isothermal_Glen.ice_softness_units = "Pascal-3 second-1";

    pism_overrides:fracture_density.constant_fd = "no";
    pism_overrides:fracture_density.constant_fd_doc = "FIXME";
    pism_overrides:fracture_density.constant_fd_option = "constant_fd";
    pism_overrides:fracture_density.constant_fd_type = "flag";

    pism_overrides:fracture_density.constant_healing = "no";
    pism_overrides:fracture_density.constant_healing_doc = "Constant healing";
    pism_overrides:fracture_density.constant_healing_option = "constant_healing";
    pism_overrides:fracture_density.constant_healing_type = "flag";

    pism_overrides:fracture_density.enabled = "no";
    pism_overrides:fracture_density.enabled_doc = "Calculation of fracture density according to stresses and strain rate field.";
    pism_overrides:fracture_density.enabled_option = "fractures";
    pism_overrides:fracture_density.enabled_type = "flag";

    pism_overrides:fracture_density.fd2d_scheme = "no";
    pism_overrides:fracture_density.fd2d_scheme_doc = "FIXME";
    pism_overrides:fracture_density.fd2d_scheme_option = "scheme_fd2d";
    pism_overrides:fracture_density.fd2d_scheme_type = "flag";

    pism_overrides:fracture_density.fracture_weighted_healing = "no";
    pism_overrides:fracture_density.fracture_weighted_healing_doc = "Fracture weighted healing";
    pism_overrides:fracture_density.fracture_weighted_healing_option = "fracture_weighted_healing";
    pism_overrides:fracture_density.fracture_weighted_healing_type = "flag";

    pism_overrides:fracture_density.include_grounded_ice = "no";
    pism_overrides:fracture_density.include_grounded_ice_doc = "model fracture density in grounded areas";
    pism_overrides:fracture_density.include_grounded_ice_option = "do_frac_on_grounded";
    pism_overrides:fracture_density.include_grounded_ice_type = "flag";

    pism_overrides:fracture_density.lefm = "no";
    pism_overrides:fracture_density.lefm_doc = "FIXME";
    pism_overrides:fracture_density.lefm_option = "lefm";
    pism_overrides:fracture_density.lefm_type = "flag";

    pism_overrides:fracture_density.max_shear_stress = "no";
    pism_overrides:fracture_density.max_shear_stress_doc = "Use the max. shear stress criterion.";
    pism_overrides:fracture_density.max_shear_stress_option = "max_shear";
    pism_overrides:fracture_density.max_shear_stress_type = "flag";

    pism_overrides:fracture_density.phi0 = 0.0;
    pism_overrides:fracture_density.phi0_doc = "FIXME";
    pism_overrides:fracture_density.phi0_option = "phi0";
    pism_overrides:fracture_density.phi0_type = "number";
    pism_overrides:fracture_density.phi0_units = "1";

    pism_overrides:fracture_density.softening_lower_limit = 1.0;
    pism_overrides:fracture_density.softening_lower_limit_doc = "epsilon in equation (6) in Albrecht and Levermann, 'Fracture-induced softening for large-scale ice dynamics'";
    pism_overrides:fracture_density.softening_lower_limit_option = "fracture_softening";
    pism_overrides:fracture_density.softening_lower_limit_type = "number";
    pism_overrides:fracture_density.softening_lower_limit_units = "1";

    pism_overrides:frontal_melt.constant.melt_rate = 1.0;
    pism_overrides:frontal_melt.constant.melt_rate_doc = "default melt rate used by the 'constant' frontal_melt model";
    pism_overrides:frontal_melt.constant.melt_rate_option = "frontal_melt_rate";
    pism_overrides:frontal_melt.constant.melt_rate_type = "number";
    pism_overrides:frontal_melt.constant.melt_rate_units = "m / day";

    pism_overrides:frontal_melt.discharge_given.file = "";
    pism_overrides:frontal_melt.discharge_given.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:frontal_melt.discharge_given.file_option = "frontal_melt_discharge_given_file";
    pism_overrides:frontal_melt.discharge_given.file_type = "string";

    pism_overrides:frontal_melt.discharge_given.period = 0;
    pism_overrides:frontal_melt.discharge_given.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:frontal_melt.discharge_given.period_option = "frontal_melt_discharge_given_period";
    pism_overrides:frontal_melt.discharge_given.period_type = "integer";
    pism_overrides:frontal_melt.discharge_given.period_units = "years";

    pism_overrides:frontal_melt.discharge_given.reference_year = 0;
    pism_overrides:frontal_melt.discharge_given.reference_year_doc = "Reference year to use when ``frontal_melt.discharge_given.period`` is active.";
    pism_overrides:frontal_melt.discharge_given.reference_year_option = "frontal_melt_discharge_given_reference_year";
    pism_overrides:frontal_melt.discharge_given.reference_year_type = "integer";
    pism_overrides:frontal_melt.discharge_given.reference_year_units = "years";

    pism_overrides:frontal_melt.given.file = "";
    pism_overrides:frontal_melt.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:frontal_melt.given.file_option = "frontal_melt_given_file";
    pism_overrides:frontal_melt.given.file_type = "string";

    pism_overrides:frontal_melt.given.period = 0;
    pism_overrides:frontal_melt.given.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:frontal_melt.given.period_option = "frontal_melt_given_period";
    pism_overrides:frontal_melt.given.period_type = "integer";
    pism_overrides:frontal_melt.given.period_units = "years";

    pism_overrides:frontal_melt.given.reference_year = 0;
    pism_overrides:frontal_melt.given.reference_year_doc = "Reference year to use when ``frontal_melt.given.period`` is active.";
    pism_overrides:frontal_melt.given.reference_year_option = "frontal_melt_given_reference_year";
    pism_overrides:frontal_melt.given.reference_year_type = "integer";
    pism_overrides:frontal_melt.given.reference_year_units = "years";

    pism_overrides:frontal_melt.include_floating_ice = "no";
    pism_overrides:frontal_melt.include_floating_ice_doc = "Apply frontal melt to all grid icy cells next to ocean cells";
    pism_overrides:frontal_melt.include_floating_ice_type = "flag";

    pism_overrides:frontal_melt.models = "";
    pism_overrides:frontal_melt.models_doc = "Comma-separated list of frontal melt models and modifiers. (Leave empty to disable.)";
    pism_overrides:frontal_melt.models_option = "frontal_melt";
    pism_overrides:frontal_melt.models_type = "string";

    pism_overrides:frontal_melt.routing.file = "";
    pism_overrides:frontal_melt.routing.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:frontal_melt.routing.file_option = "frontal_melt_routing_file";
    pism_overrides:frontal_melt.routing.file_type = "string";

    pism_overrides:frontal_melt.routing.parameter_a = 3e-4;
    pism_overrides:frontal_melt.routing.parameter_a_doc = "parameter A in eqn. 1 in :cite:`Xu2013`";
    pism_overrides:frontal_melt.routing.parameter_a_type = "number";
    pism_overrides:frontal_melt.routing.parameter_a_units = "m-alpha day^(alpha-1) Celsius-beta";

    pism_overrides:frontal_melt.routing.parameter_b = 0.15;
    pism_overrides:frontal_melt.routing.parameter_b_doc = "parameter B in eqn. 1 in :cite:`Xu2013`";
    pism_overrides:frontal_melt.routing.parameter_b_type = "number";
    pism_overrides:frontal_melt.routing.parameter_b_units = "m day^(alpha-1) Celsius-beta";

    pism_overrides:frontal_melt.routing.period = 0;
    pism_overrides:frontal_melt.routing.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:frontal_melt.routing.period_option = "frontal_melt_routing_period";
    pism_overrides:frontal_melt.routing.period_type = "integer";
    pism_overrides:frontal_melt.routing.period_units = "years";

    pism_overrides:frontal_melt.routing.power_alpha = 0.39;
    pism_overrides:frontal_melt.routing.power_alpha_doc = "exponent `\\alpha` in eqn. 1 in :cite:`Xu2013`";
    pism_overrides:frontal_melt.routing.power_alpha_type = "number";
    pism_overrides:frontal_melt.routing.power_alpha_units = "1";

    pism_overrides:frontal_melt.routing.power_beta = 1.18;
    pism_overrides:frontal_melt.routing.power_beta_doc = "exponent `\\beta` in eqn. 1 in :cite:`Xu2013`";
    pism_overrides:frontal_melt.routing.power_beta_type = "number";
    pism_overrides:frontal_melt.routing.power_beta_units = "1";

    pism_overrides:frontal_melt.routing.reference_year = 0;
    pism_overrides:frontal_melt.routing.reference_year_doc = "Reference year to use when ``frontal_melt.routing.period`` is active.";
    pism_overrides:frontal_melt.routing.reference_year_option = "frontal_melt_routing_reference_year";
    pism_overrides:frontal_melt.routing.reference_year_type = "integer";
    pism_overrides:frontal_melt.routing.reference_year_units = "years";

    pism_overrides:geometry.front_retreat.prescribed.file = "";
    pism_overrides:geometry.front_retreat.prescribed.file_doc = "Name of the file containing the maximum ice extent mask `land_ice_area_fraction_retreat`";
    pism_overrides:geometry.front_retreat.prescribed.file_option = "front_retreat_file";
    pism_overrides:geometry.front_retreat.prescribed.file_type = "string";

    pism_overrides:geometry.front_retreat.prescribed.period = 0;
    pism_overrides:geometry.front_retreat.prescribed.period_doc = "Length of the period of the front retreat data. Set to zero to disable.";
    pism_overrides:geometry.front_retreat.prescribed.period_type = "integer";
    pism_overrides:geometry.front_retreat.prescribed.period_units = "years";

    pism_overrides:geometry.front_retreat.prescribed.reference_year = 0;
    pism_overrides:geometry.front_retreat.prescribed.reference_year_doc = "Reference year to use when `geometry.front_retreat.prescribed.period` is active.";
    pism_overrides:geometry.front_retreat.prescribed.reference_year_type = "integer";
    pism_overrides:geometry.front_retreat.prescribed.reference_year_units = "years";

    pism_overrides:geometry.front_retreat.use_cfl = "false";
    pism_overrides:geometry.front_retreat.use_cfl_doc = "apply CFL criterion for eigen-calving rate front retreat";
    pism_overrides:geometry.front_retreat.use_cfl_option = "front_retreat_cfl";
    pism_overrides:geometry.front_retreat.use_cfl_type = "flag";

    pism_overrides:geometry.front_retreat.wrap_around = "false";
    pism_overrides:geometry.front_retreat.wrap_around_doc = "If true, wrap around domain boundaries. This may be needed in some regional synthetic geometry setups.";
    pism_overrides:geometry.front_retreat.wrap_around_option = "front_retreat_wrap_around";
    pism_overrides:geometry.front_retreat.wrap_around_type = "flag";

    pism_overrides:geometry.grounded_cell_fraction  = "false";
    pism_overrides:geometry.grounded_cell_fraction_doc = "Linear interpolation scheme ('LI' in Gladstone et al. 2010) expanded to two dimensions is used if switched on in order to evaluate the position of the grounding line on a subgrid scale.";
    pism_overrides:geometry.grounded_cell_fraction_option = "subgl";
    pism_overrides:geometry.grounded_cell_fraction_type = "flag";

    pism_overrides:geometry.ice_free_thickness_standard = 0.01;
    pism_overrides:geometry.ice_free_thickness_standard_doc = "If ice is thinner than this standard then the mask is set to MASK_ICE_FREE_BEDROCK or MASK_ICE_FREE_OCEAN.";
    pism_overrides:geometry.ice_free_thickness_standard_type = "number";
    pism_overrides:geometry.ice_free_thickness_standard_units = "meters";

    pism_overrides:geometry.part_grid.enabled = "no";
    pism_overrides:geometry.part_grid.enabled_doc = "apply partially filled grid cell scheme";
    pism_overrides:geometry.part_grid.enabled_option = "part_grid";
    pism_overrides:geometry.part_grid.enabled_type = "flag";

    pism_overrides:geometry.part_grid.max_iterations = 10;
    pism_overrides:geometry.part_grid.max_iterations_doc = "maximum number of residual redistribution iterations";
    pism_overrides:geometry.part_grid.max_iterations_type = "integer";
    pism_overrides:geometry.part_grid.max_iterations_units = "count";

    pism_overrides:geometry.remove_icebergs = "no";
    pism_overrides:geometry.remove_icebergs_doc = "identify and kill detached ice-shelf areas";
    pism_overrides:geometry.remove_icebergs_option = "kill_icebergs";
    pism_overrides:geometry.remove_icebergs_type = "flag";

    pism_overrides:geometry.update.enabled = "yes";
    pism_overrides:geometry.update.enabled_doc = "Solve the mass conservation equation";
    pism_overrides:geometry.update.enabled_option = "mass";
    pism_overrides:geometry.update.enabled_type = "flag";

    pism_overrides:geometry.update.use_basal_melt_rate = "yes";
    pism_overrides:geometry.update.use_basal_melt_rate_doc = "Include basal melt rate in the continuity equation";
    pism_overrides:geometry.update.use_basal_melt_rate_option = "bmr_in_cont";
    pism_overrides:geometry.update.use_basal_melt_rate_type = "flag";

    pism_overrides:grid.Lbz = 1000;
    pism_overrides:grid.Lbz_doc = "Thickness of the thermal bedrock layer. (Inactive if ``grid.Mbz`` < 2)";
    pism_overrides:grid.Lbz_option = "Lbz";
    pism_overrides:grid.Lbz_type = "number";
    pism_overrides:grid.Lbz_units = "meters";

    pism_overrides:grid.Lx = 1500e3;
    pism_overrides:grid.Lx_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_overrides:grid.Lx_type = "number";
    pism_overrides:grid.Lx_units = "meters";

    pism_overrides:grid.Ly = 1500e3;
    pism_overrides:grid.Ly_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_overrides:grid.Ly_type = "number";
    pism_overrides:grid.Ly_units = "meters";

    pism_overrides:grid.Lz = 4000;
    pism_overrides:grid.Lz_doc = "Height of the computational domain.";
    pism_overrides:grid.Lz_option = "Lz";
    pism_overrides:grid.Lz_type = "number";
    pism_overrides:grid.Lz_units = "meters";

    pism_overrides:grid.Mbz = 1;
    pism_overrides:grid.Mbz_doc = "Number of thermal bedrock layers; 1 level corresponds to no bedrock.";
    pism_overrides:grid.Mbz_option = "Mbz";
    pism_overrides:grid.Mbz_type = "integer";
    pism_overrides:grid.Mbz_units = "count";

    pism_overrides:grid.Mx = 61;
    pism_overrides:grid.Mx_doc = "Number of grid points in the x direction.";
    pism_overrides:grid.Mx_option = "Mx";
    pism_overrides:grid.Mx_type = "integer";
    pism_overrides:grid.Mx_units = "count";

    pism_overrides:grid.My = 61;
    pism_overrides:grid.My_doc = "Number of grid points in the y direction.";
    pism_overrides:grid.My_option = "My";
    pism_overrides:grid.My_type = "integer";
    pism_overrides:grid.My_units = "count";

    pism_overrides:grid.Mz = 31;
    pism_overrides:grid.Mz_doc = "Number of vertical grid levels in the ice.";
    pism_overrides:grid.Mz_option = "Mz";
    pism_overrides:grid.Mz_type = "integer";
    pism_overrides:grid.Mz_units = "count";

    pism_overrides:grid.allow_extrapolation = "no";
    pism_overrides:grid.allow_extrapolation_doc = "Allow extrapolation during regridding.";
    pism_overrides:grid.allow_extrapolation_option = "allow_extrapolation";
    pism_overrides:grid.allow_extrapolation_type = "flag";

    pism_overrides:grid.ice_vertical_spacing = "quadratic";
    pism_overrides:grid.ice_vertical_spacing_choices = "quadratic,equal";
    pism_overrides:grid.ice_vertical_spacing_doc = "vertical spacing in the ice";
    pism_overrides:grid.ice_vertical_spacing_option = "z_spacing";
    pism_overrides:grid.ice_vertical_spacing_type = "keyword";

    pism_overrides:grid.lambda = 4.0;
    pism_overrides:grid.lambda_doc = "Vertical grid spacing parameter. Roughly equal to the factor by which the grid is coarser at an end away from the ice-bedrock interface.";
    pism_overrides:grid.lambda_type = "number";
    pism_overrides:grid.lambda_units = "pure number";

    pism_overrides:grid.max_stencil_width = 2;
    pism_overrides:grid.max_stencil_width_doc = "Maximum width of the finite-difference stencil used in PISM.";
    pism_overrides:grid.max_stencil_width_type = "integer";
    pism_overrides:grid.max_stencil_width_units = "count";

    pism_overrides:grid.periodicity = "xy";
    pism_overrides:grid.periodicity_choices = "none,x,y,xy";
    pism_overrides:grid.periodicity_doc = "horizontal grid periodicity";
    pism_overrides:grid.periodicity_option = "periodicity";
    pism_overrides:grid.periodicity_type = "keyword";

    pism_overrides:grid.recompute_longitude_and_latitude = "yes";
    pism_overrides:grid.recompute_longitude_and_latitude_doc = "Re-compute longitude and latitude using grid information and provided projection parameters. Requires PROJ.";
    pism_overrides:grid.recompute_longitude_and_latitude_type = "flag";

    pism_overrides:grid.registration = "center";
    pism_overrides:grid.registration_choices = "center,corner";
    pism_overrides:grid.registration_doc = "horizontal grid registration";
    pism_overrides:grid.registration_type = "keyword";

    pism_overrides:hydrology.add_water_input_to_till_storage = "yes";
    pism_overrides:hydrology.add_water_input_to_till_storage_doc = "Add surface input to water stored in till. If no it will be added to the transportable water.";
    pism_overrides:hydrology.add_water_input_to_till_storage_type = "flag";

    pism_overrides:hydrology.cavitation_opening_coefficient = 0.5;
    pism_overrides:hydrology.cavitation_opening_coefficient_doc = "c_1 in notes; coefficient of cavitation opening term in evolution of layer thickness in hydrology::Distributed";
    pism_overrides:hydrology.cavitation_opening_coefficient_option = "hydrology_cavitation_opening_coefficient";
    pism_overrides:hydrology.cavitation_opening_coefficient_type = "number";
    pism_overrides:hydrology.cavitation_opening_coefficient_units = "meter-1";

    pism_overrides:hydrology.creep_closure_coefficient = 0.04;
    pism_overrides:hydrology.creep_closure_coefficient_doc = "c_2 in notes; coefficient of creep closure term in evolution of layer thickness in hydrology::Distributed";
    pism_overrides:hydrology.creep_closure_coefficient_option = "hydrology_creep_closure_coefficient";
    pism_overrides:hydrology.creep_closure_coefficient_type = "number";
    pism_overrides:hydrology.creep_closure_coefficient_units = "pure number";

    pism_overrides:hydrology.distributed.init_p_from_steady = "no";
    pism_overrides:hydrology.distributed.init_p_from_steady_doc = "if 'yes', initialize subglacial water pressure from P(W) formula that applies in steady state";
    pism_overrides:hydrology.distributed.init_p_from_steady_option = "hydrology_init_p_form_steady";
    pism_overrides:hydrology.distributed.init_p_from_steady_type = "flag";

    pism_overrides:hydrology.distributed.sliding_speed_file = "";
    pism_overrides:hydrology.distributed.sliding_speed_file_doc = "name of the file containing velbase_mag, the basal sliding speed to use with :literal:`hydrology.distributed.init_p_from_steady`";
    pism_overrides:hydrology.distributed.sliding_speed_file_option = "hydrology_sliding_speed_file";
    pism_overrides:hydrology.distributed.sliding_speed_file_type = "string";

    pism_overrides:hydrology.gradient_power_in_flux = 1.5;
    pism_overrides:hydrology.gradient_power_in_flux_doc = "power `\\beta` in Darcy's law `q = - k W^{\\alpha} |\\nabla \\psi|^{\\beta-2} \\nabla \\psi`, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_overrides:hydrology.gradient_power_in_flux_option = "hydrology_gradient_power_in_flux";
    pism_overrides:hydrology.gradient_power_in_flux_type = "number";
    pism_overrides:hydrology.gradient_power_in_flux_units = "pure number";

    pism_overrides:hydrology.hydraulic_conductivity = 0.001;
    pism_overrides:hydrology.hydraulic_conductivity_doc = "= k in notes; lateral conductivity, in Darcy's law, for subglacial water layer; units depend on powers alpha = hydrology.thickness_power_in_flux and beta = hydrology_potential_gradient_power_in_flux; used by hydrology::Routing and hydrology::Distributed";
    pism_overrides:hydrology.hydraulic_conductivity_option = "hydrology_hydraulic_conductivity";
    pism_overrides:hydrology.hydraulic_conductivity_type = "number";
    pism_overrides:hydrology.hydraulic_conductivity_units = "`m^{2 \\beta - \\alpha} s^{2 \\beta - 3} kg^{1-\\beta}`";

    pism_overrides:hydrology.maximum_time_step = 1.0;
    pism_overrides:hydrology.maximum_time_step_doc = "maximum allowed time step length used by hydrology::Routing and hydrology::Distributed";
    pism_overrides:hydrology.maximum_time_step_type = "number";
    pism_overrides:hydrology.maximum_time_step_units = "years";

    pism_overrides:hydrology.model = "null";
    pism_overrides:hydrology.model_choices = "null,routing,steady,distributed";
    pism_overrides:hydrology.model_doc = "Basal hydrology sub-model.";
    pism_overrides:hydrology.model_option = "hydrology";
    pism_overrides:hydrology.model_type = "keyword";

    pism_overrides:hydrology.null_diffuse_till_water = "no";
    pism_overrides:hydrology.null_diffuse_till_water_doc = "Diffuse stored till water laterally. See equation (11) of :cite:`BBssasliding`";
    pism_overrides:hydrology.null_diffuse_till_water_type = "flag";

    pism_overrides:hydrology.null_diffusion_distance = 2e4;
    pism_overrides:hydrology.null_diffusion_distance_doc = "diffusion distance for till water thickness; see equation (11) in :cite:`BBssasliding`; only active if hydrology.null_diffuse_till_water is set";
    pism_overrides:hydrology.null_diffusion_distance_type = "number";
    pism_overrides:hydrology.null_diffusion_distance_units = "meters";

    pism_overrides:hydrology.null_diffusion_time = 1000.0;
    pism_overrides:hydrology.null_diffusion_time_doc = "diffusion time for till water thickness; see equation (11) in :cite:`BBssasliding`; only active if hydrology.null_diffuse_till_water is set";
    pism_overrides:hydrology.null_diffusion_time_type = "number";
    pism_overrides:hydrology.null_diffusion_time_units = "years";

    pism_overrides:hydrology.null_strip_width = -1.0;
    pism_overrides:hydrology.null_strip_width_doc = "if negative then mechanism is inactive; width of strip around computational domain in which water velocity and water amount are set to zero; used by hydrology::Routing and hydrology::Distributed";
    pism_overrides:hydrology.null_strip_width_type = "number";
    pism_overrides:hydrology.null_strip_width_units = "meters";

    pism_overrides:hydrology.regularizing_porosity = 0.01;
    pism_overrides:hydrology.regularizing_porosity_doc = "phi_0 in notes; regularizes pressure equation by multiplying time derivative term";
    pism_overrides:hydrology.regularizing_porosity_option = "hydrology_regularizing_porosity";
    pism_overrides:hydrology.regularizing_porosity_type = "number";
    pism_overrides:hydrology.regularizing_porosity_units = "pure number";

    pism_overrides:hydrology.roughness_scale = 0.1;
    pism_overrides:hydrology.roughness_scale_doc = "W_r in notes; roughness scale determining maximum amount of cavitation opening in hydrology::Distributed";
    pism_overrides:hydrology.roughness_scale_option = "hydrology_roughness_scale";
    pism_overrides:hydrology.roughness_scale_type = "number";
    pism_overrides:hydrology.roughness_scale_units = "meters";

    pism_overrides:hydrology.routing.include_floating_ice = "no";
    pism_overrides:hydrology.routing.include_floating_ice_doc = "Route subglacial water under ice shelves. This may be appropriate if a shelf is close to floatation. Note that this has no effect on ice flow.";
    pism_overrides:hydrology.routing.include_floating_ice_type = "flag";

    pism_overrides:hydrology.steady.flux_update_interval = 1.0;
    pism_overrides:hydrology.steady.flux_update_interval_doc = "interval between updates of the steady state flux";
    pism_overrides:hydrology.steady.flux_update_interval_type = "number";
    pism_overrides:hydrology.steady.flux_update_interval_units = "years";

    pism_overrides:hydrology.steady.input_rate_scaling = 1e7;
    pism_overrides:hydrology.steady.input_rate_scaling_doc = "input rate scaling";
    pism_overrides:hydrology.steady.input_rate_scaling_type = "number";
    pism_overrides:hydrology.steady.input_rate_scaling_units = "seconds";

    pism_overrides:hydrology.steady.n_iterations = 7500;
    pism_overrides:hydrology.steady.n_iterations_doc = "maxinum number of iterations to use in while estimating steady-state water flux";
    pism_overrides:hydrology.steady.n_iterations_type = "integer";
    pism_overrides:hydrology.steady.n_iterations_units = "count";

    pism_overrides:hydrology.steady.potential_delta = 10000.0;
    pism_overrides:hydrology.steady.potential_delta_doc = "potential adjustment used to fill sinks (smaller values require more iterations but produce fewer artifacts)";
    pism_overrides:hydrology.steady.potential_delta_type = "number";
    pism_overrides:hydrology.steady.potential_delta_units = "Pa";

    pism_overrides:hydrology.steady.potential_n_iterations = 1000;
    pism_overrides:hydrology.steady.potential_n_iterations_doc = "maxinum number of iterations to take while pre-processing hydraulic potential";
    pism_overrides:hydrology.steady.potential_n_iterations_type = "integer";
    pism_overrides:hydrology.steady.potential_n_iterations_units = "count";

    pism_overrides:hydrology.steady.volume_ratio = 0.1;
    pism_overrides:hydrology.steady.volume_ratio_doc = "water volume ratio used as the stopping criterion";
    pism_overrides:hydrology.steady.volume_ratio_type = "number";
    pism_overrides:hydrology.steady.volume_ratio_units = "1";

    pism_overrides:hydrology.surface_input.file = "";
    pism_overrides:hydrology.surface_input.file_doc = "Name of the file containing ``water_input_rate``, the rate at which water from the ice surface is added to the subglacial hydrology system";
    pism_overrides:hydrology.surface_input.file_type = "string";

    pism_overrides:hydrology.surface_input.period = 0;
    pism_overrides:hydrology.surface_input.period_doc = "Length of the period of the water input rate. Set to zero to disable.";
    pism_overrides:hydrology.surface_input.period_type = "integer";
    pism_overrides:hydrology.surface_input.period_units = "years";

    pism_overrides:hydrology.surface_input.reference_year = 0;
    pism_overrides:hydrology.surface_input.reference_year_doc = "Reference year to use when ``hydrology.surface_input.period`` is active.";
    pism_overrides:hydrology.surface_input.reference_year_type = "integer";
    pism_overrides:hydrology.surface_input.reference_year_units = "years";

    pism_overrides:hydrology.surface_input_from_runoff = "no";
    pism_overrides:hydrology.surface_input_from_runoff_doc = "Use surface runoff as surface input.";
    pism_overrides:hydrology.surface_input_from_runoff_type = "flag";

    pism_overrides:hydrology.thickness_power_in_flux = 1.25;
    pism_overrides:hydrology.thickness_power_in_flux_doc = "power `\\alpha` in Darcy's law `q = - k W^{\\alpha} |\\nabla \\psi|^{\\beta-2} \\nabla \\psi`, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_overrides:hydrology.thickness_power_in_flux_option = "hydrology_thickness_power_in_flux";
    pism_overrides:hydrology.thickness_power_in_flux_type = "number";
    pism_overrides:hydrology.thickness_power_in_flux_units = "1";

    pism_overrides:hydrology.tillwat_decay_rate = 1.0;
    pism_overrides:hydrology.tillwat_decay_rate_doc = "rate at which tillwat is reduced to zero, in absence of other effects like input";
    pism_overrides:hydrology.tillwat_decay_rate_option = "hydrology_tillwat_decay_rate";
    pism_overrides:hydrology.tillwat_decay_rate_type = "number";
    pism_overrides:hydrology.tillwat_decay_rate_units = "mm / year";

    pism_overrides:hydrology.tillwat_max = 2.0;
    pism_overrides:hydrology.tillwat_max_doc = "maximum effective thickness of the water stored in till";
    pism_overrides:hydrology.tillwat_max_option = "hydrology_tillwat_max";
    pism_overrides:hydrology.tillwat_max_type = "number";
    pism_overrides:hydrology.tillwat_max_units = "meters";

    pism_overrides:hydrology.use_const_bmelt = "no";
    pism_overrides:hydrology.use_const_bmelt_doc = "if 'yes', subglacial hydrology model sees basal melt rate which is constant and given by hydrology.const_bmelt";
    pism_overrides:hydrology.use_const_bmelt_option = "hydrology_use_const_bmelt";
    pism_overrides:hydrology.use_const_bmelt_type = "flag";

    pism_overrides:input.bootstrap = "no";
    pism_overrides:input.bootstrap_doc = "It true, use bootstrapping heuristics when initializing PISM.";
    pism_overrides:input.bootstrap_option = "bootstrap";
    pism_overrides:input.bootstrap_type = "flag";

    pism_overrides:input.file = "";
    pism_overrides:input.file_doc = "Input file name";
    pism_overrides:input.file_option = "i";
    pism_overrides:input.file_type = "string";

    pism_overrides:input.forcing.buffer_size = 60;
    pism_overrides:input.forcing.buffer_size_doc = "number of 2D climate forcing records to keep in memory; = 5 years of monthly records";
    pism_overrides:input.forcing.buffer_size_type = "integer";
    pism_overrides:input.forcing.buffer_size_units = "count";

    pism_overrides:input.forcing.evaluations_per_year = 52;
    pism_overrides:input.forcing.evaluations_per_year_doc = "length of the time-series used to compute temporal averages of forcing data (such as mean annual temperature)";
    pism_overrides:input.forcing.evaluations_per_year_type = "integer";
    pism_overrides:input.forcing.evaluations_per_year_units = "count";

    pism_overrides:input.regrid.file = "";
    pism_overrides:input.regrid.file_doc = "Regridding (input) file name";
    pism_overrides:input.regrid.file_option = "regrid_file";
    pism_overrides:input.regrid.file_type = "string";

    pism_overrides:input.regrid.vars = "";
    pism_overrides:input.regrid.vars_doc = "Comma-separated list of variables to regrid. Leave empty to regrid all model state variables.";
    pism_overrides:input.regrid.vars_option = "regrid_vars";
    pism_overrides:input.regrid.vars_type = "string";

    pism_overrides:inverse.design.cH1     = 0;
    pism_overrides:inverse.design.cH1_doc = "weight of derivative part of an H1 norm for inversion design variables";
    pism_overrides:inverse.design.cH1_option = "inv_design_cH1";
    pism_overrides:inverse.design.cH1_type = "number";
    pism_overrides:inverse.design.cH1_units = "1";

    pism_overrides:inverse.design.cL2 = 1;
    pism_overrides:inverse.design.cL2_doc = "weight of derivative-free part of an H1 norm for inversion design variables";
    pism_overrides:inverse.design.cL2_option = "inv_design_cL2";
    pism_overrides:inverse.design.cL2_type = "number";
    pism_overrides:inverse.design.cL2_units = "1";

    pism_overrides:inverse.design.func = "sobolevH1";
    pism_overrides:inverse.design.func_choices = "sobolevH1,tv";
    pism_overrides:inverse.design.func_doc = "functional used for inversion design variables";
    pism_overrides:inverse.design.func_option = "inv_design_func";
    pism_overrides:inverse.design.func_type = "keyword";

    pism_overrides:inverse.design.param = "exp";
    pism_overrides:inverse.design.param_choices = "ident,trunc,square,exp";
    pism_overrides:inverse.design.param_doc = "parameterization of design variables used during inversion";
    pism_overrides:inverse.design.param_option = "inv_design_param";
    pism_overrides:inverse.design.param_type = "keyword";

    pism_overrides:inverse.design.param_hardav_eps = 1e4;
    pism_overrides:inverse.design.param_hardav_eps_doc = "tiny vertically-averaged hardness used as a substitute for 0 in some tauc parameterizations";
    pism_overrides:inverse.design.param_hardav_eps_type = "number";
    pism_overrides:inverse.design.param_hardav_eps_units = "Pascal second^(1/3)";

    pism_overrides:inverse.design.param_hardav_scale = 1e8;
    pism_overrides:inverse.design.param_hardav_scale_doc = "typical size of ice hardness";
    pism_overrides:inverse.design.param_hardav_scale_type = "number";
    pism_overrides:inverse.design.param_hardav_scale_units = "Pascal second^(1/3)";

    pism_overrides:inverse.design.param_tauc_eps = 100;
    pism_overrides:inverse.design.param_tauc_eps_doc = "tiny yield stress used as a substitute for 0 in some tauc parameterizations";
    pism_overrides:inverse.design.param_tauc_eps_type = "number";
    pism_overrides:inverse.design.param_tauc_eps_units = "Pascal";

    pism_overrides:inverse.design.param_tauc_scale = 100000;
    pism_overrides:inverse.design.param_tauc_scale_doc = "typical size of yield stresses";
    pism_overrides:inverse.design.param_tauc_scale_type = "number";
    pism_overrides:inverse.design.param_tauc_scale_units = "Pascal";

    pism_overrides:inverse.design.param_trunc_hardav0 = 1e6;
    pism_overrides:inverse.design.param_trunc_hardav0_doc = "transition point of change to linear behaviour for design variable parameterization type 'trunc'";
    pism_overrides:inverse.design.param_trunc_hardav0_type = "number";
    pism_overrides:inverse.design.param_trunc_hardav0_units = "Pascal second^(1/3)";

    pism_overrides:inverse.design.param_trunc_tauc0 = 1000;
    pism_overrides:inverse.design.param_trunc_tauc0_doc = "transition point of change to linear behaviour for design variable parameterization type 'trunc'";
    pism_overrides:inverse.design.param_trunc_tauc0_type = "number";
    pism_overrides:inverse.design.param_trunc_tauc0_units = "Pascal";

    pism_overrides:inverse.log_ratio_scale = 10;
    pism_overrides:inverse.log_ratio_scale_doc = "Reference scale for log-ratio functionals";
    pism_overrides:inverse.log_ratio_scale_option = "inv_log_ratio_scale";
    pism_overrides:inverse.log_ratio_scale_type = "number";
    pism_overrides:inverse.log_ratio_scale_units = "pure number";

    pism_overrides:inverse.max_iterations = 1000;
    pism_overrides:inverse.max_iterations_doc = "maximum iteration count";
    pism_overrides:inverse.max_iterations_option = "inv_max_it";
    pism_overrides:inverse.max_iterations_type = "integer";
    pism_overrides:inverse.max_iterations_units = "count";

    pism_overrides:inverse.ssa.hardav_max = 1e10;
    pism_overrides:inverse.ssa.hardav_max_doc = "Maximum allowed value of hardav for inversions with bound constraints";
    pism_overrides:inverse.ssa.hardav_max_type = "number";
    pism_overrides:inverse.ssa.hardav_max_units = "Pascal second^(1/3)";

    pism_overrides:inverse.ssa.hardav_min = 0;
    pism_overrides:inverse.ssa.hardav_min_doc = "Minimum allowed value of hardav for inversions with bound constraints";
    pism_overrides:inverse.ssa.hardav_min_type = "number";
    pism_overrides:inverse.ssa.hardav_min_units = "Pascal second^(1/3)";

    pism_overrides:inverse.ssa.length_scale = 50e3;
    pism_overrides:inverse.ssa.length_scale_doc = "typical length scale for rescaling derivative norms";
    pism_overrides:inverse.ssa.length_scale_type = "number";
    pism_overrides:inverse.ssa.length_scale_units = "meters";

    pism_overrides:inverse.ssa.method = "tikhonov_lmvm";
    pism_overrides:inverse.ssa.method_choices = "sd,nlcg,ign,tikhonov_lmvm,tikhonov_cg,tikhonov_blmvm,tikhonov_lcl,tikhonov_gn";
    pism_overrides:inverse.ssa.method_doc = "algorithm to use for SSA inversions";
    pism_overrides:inverse.ssa.method_option = "inv_method";
    pism_overrides:inverse.ssa.method_type = "keyword";

    pism_overrides:inverse.ssa.tauc_max = 5e7;
    pism_overrides:inverse.ssa.tauc_max_doc = "Maximum allowed value of tauc for inversions with bound constraints";
    pism_overrides:inverse.ssa.tauc_max_type = "number";
    pism_overrides:inverse.ssa.tauc_max_units = "Pascal";

    pism_overrides:inverse.ssa.tauc_min = 0;
    pism_overrides:inverse.ssa.tauc_min_doc = "Minimum allowed value of tauc for inversions with bound constraints";
    pism_overrides:inverse.ssa.tauc_min_type = "number";
    pism_overrides:inverse.ssa.tauc_min_units = "Pascal";

    pism_overrides:inverse.ssa.tv_exponent = 1.2;
    pism_overrides:inverse.ssa.tv_exponent_doc = "Lebesgue exponent for pseudo-TV norm";
    pism_overrides:inverse.ssa.tv_exponent_option = "inv_ssa_tv_exponent";
    pism_overrides:inverse.ssa.tv_exponent_type = "number";
    pism_overrides:inverse.ssa.tv_exponent_units = "pure number";

    pism_overrides:inverse.ssa.velocity_eps = 0.1;
    pism_overrides:inverse.ssa.velocity_eps_doc = "tiny size of ice velocities during inversion";
    pism_overrides:inverse.ssa.velocity_eps_type = "number";
    pism_overrides:inverse.ssa.velocity_eps_units = "meter / year";

    pism_overrides:inverse.ssa.velocity_scale = 100;
    pism_overrides:inverse.ssa.velocity_scale_doc = "typical size of ice velocities expected during inversion";
    pism_overrides:inverse.ssa.velocity_scale_type = "number";
    pism_overrides:inverse.ssa.velocity_scale_units = "meter / year";

    pism_overrides:inverse.state_func = "meansquare";
    pism_overrides:inverse.state_func_choices = "meansquare,log_ratio,log_relative";
    pism_overrides:inverse.state_func_doc = "functional used for inversion design variables";
    pism_overrides:inverse.state_func_option = "inv_state_func";
    pism_overrides:inverse.state_func_type = "keyword";

    pism_overrides:inverse.target_misfit = 100;
    pism_overrides:inverse.target_misfit_doc = "desired root misfit for SSA inversions";
    pism_overrides:inverse.target_misfit_option = "inv_target_misfit";
    pism_overrides:inverse.target_misfit_type = "number";
    pism_overrides:inverse.target_misfit_units = "meter / year";

    pism_overrides:inverse.tikhonov.atol = 1e-10;
    pism_overrides:inverse.tikhonov.atol_doc = "absolute threshold for Tikhonov stopping criterion";
    pism_overrides:inverse.tikhonov.atol_option = "tikhonov_atol";
    pism_overrides:inverse.tikhonov.atol_type = "number";
    pism_overrides:inverse.tikhonov.atol_units = "meter / year";

    pism_overrides:inverse.tikhonov.penalty_weight = 1;
    pism_overrides:inverse.tikhonov.penalty_weight_doc = "penalty parameter for Tikhonov inversion";
    pism_overrides:inverse.tikhonov.penalty_weight_option = "tikhonov_penalty";
    pism_overrides:inverse.tikhonov.penalty_weight_type = "number";
    pism_overrides:inverse.tikhonov.penalty_weight_units = "1";

    pism_overrides:inverse.tikhonov.ptol = 0.1;
    pism_overrides:inverse.tikhonov.ptol_doc = "threshold for reaching desired misfit for adaptive Tikhonov algorithms";
    pism_overrides:inverse.tikhonov.ptol_option = "tikhonov_ptol";
    pism_overrides:inverse.tikhonov.ptol_type = "number";
    pism_overrides:inverse.tikhonov.ptol_units = "pure number";

    pism_overrides:inverse.tikhonov.rtol = 5e-2;
    pism_overrides:inverse.tikhonov.rtol_doc = "relative threshold for Tikhonov stopping criterion";
    pism_overrides:inverse.tikhonov.rtol_option = "tikhonov_rtol";
    pism_overrides:inverse.tikhonov.rtol_type = "number";
    pism_overrides:inverse.tikhonov.rtol_units = "1";

    pism_overrides:inverse.use_design_prior = "yes";
    pism_overrides:inverse.use_design_prior_doc = "Use prior from inverse data file as initial guess.";
    pism_overrides:inverse.use_design_prior_option = "inv_use_design_prior";
    pism_overrides:inverse.use_design_prior_type = "flag";

    pism_overrides:inverse.use_zeta_fixed_mask = "yes";
    pism_overrides:inverse.use_zeta_fixed_mask_doc = "Enforce locations where the parameterized design variable should be fixed. (Automatically determined if not provided)";
    pism_overrides:inverse.use_zeta_fixed_mask_option = "inv_use_zeta_fixed_mask";
    pism_overrides:inverse.use_zeta_fixed_mask_type = "flag";

    pism_overrides:ocean.always_grounded = "no";
    pism_overrides:ocean.always_grounded_doc = "Dry (ocean-less) simulation; ice is considered grounded regardless of ice thickness, bed elevation, and sea level.";
    pism_overrides:ocean.always_grounded_option = "dry";
    pism_overrides:ocean.always_grounded_type = "flag";

    pism_overrides:ocean.anomaly.file = "";
    pism_overrides:ocean.anomaly.file_doc = "Name of the file containing shelf basal mass flux offset fields.";
    pism_overrides:ocean.anomaly.file_option = "ocean_anomaly_file";
    pism_overrides:ocean.anomaly.file_type = "string";

    pism_overrides:ocean.anomaly.period = 0;
    pism_overrides:ocean.anomaly.period_doc = "Length of the period of the ocean forcing data. Set to zero to disable.";
    pism_overrides:ocean.anomaly.period_option = "ocean_anomaly_period";
    pism_overrides:ocean.anomaly.period_type = "integer";
    pism_overrides:ocean.anomaly.period_units = "years";

    pism_overrides:ocean.anomaly.reference_year = 0;
    pism_overrides:ocean.anomaly.reference_year_doc = "Reference year to use when ``ocean.anomaly.period`` is active.";
    pism_overrides:ocean.anomaly.reference_year_option = "ocean_anomaly_reference_year";
    pism_overrides:ocean.anomaly.reference_year_type = "integer";
    pism_overrides:ocean.anomaly.reference_year_units = "years";

    pism_overrides:ocean.cache.update_interval = 10;
    pism_overrides:ocean.cache.update_interval_doc = "update interval of the 'cache' ocean modifier";
    pism_overrides:ocean.cache.update_interval_option = "ocean_cache_update_interval";
    pism_overrides:ocean.cache.update_interval_type = "integer";
    pism_overrides:ocean.cache.update_interval_units = "years";

    pism_overrides:ocean.constant.melange_back_pressure_fraction = 0.0;
    pism_overrides:ocean.constant.melange_back_pressure_fraction_doc = "default melange back pressure fraction in the 'contant' ocean model";
    pism_overrides:ocean.constant.melange_back_pressure_fraction_type = "number";
    pism_overrides:ocean.constant.melange_back_pressure_fraction_units = "1";

    pism_overrides:ocean.constant.melt_rate = 0.05191419359084029;
    pism_overrides:ocean.constant.melt_rate_doc = "default melt rate used by the 'constant' ocean model (computed as `Q / (L \\rho_i)`)";
    pism_overrides:ocean.constant.melt_rate_option = "shelf_base_melt_rate";
    pism_overrides:ocean.constant.melt_rate_type = "number";
    pism_overrides:ocean.constant.melt_rate_units = "m / year";

    pism_overrides:ocean.delta_T.file = "";
    pism_overrides:ocean.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_overrides:ocean.delta_T.file_option = "ocean_delta_T_file";
    pism_overrides:ocean.delta_T.file_type = "string";

    pism_overrides:ocean.delta_T.period = 0;
    pism_overrides:ocean.delta_T.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.delta_T.period_option = "ocean_delta_T_period";
    pism_overrides:ocean.delta_T.period_type = "integer";
    pism_overrides:ocean.delta_T.period_units = "years";

    pism_overrides:ocean.delta_T.reference_year = 0;
    pism_overrides:ocean.delta_T.reference_year_doc = "Reference year to use when ``ocean.delta_T.period`` is active.";
    pism_overrides:ocean.delta_T.reference_year_option = "ocean_delta_T_reference_year";
    pism_overrides:ocean.delta_T.reference_year_type = "integer";
    pism_overrides:ocean.delta_T.reference_year_units = "years";

    pism_overrides:ocean.delta_mass_flux.file = "";
    pism_overrides:ocean.delta_mass_flux.file_doc = "Name of the file containing sub-shelf mass flux offsets.";
    pism_overrides:ocean.delta_mass_flux.file_option = "ocean_delta_mass_flux_file";
    pism_overrides:ocean.delta_mass_flux.file_type = "string";

    pism_overrides:ocean.delta_mass_flux.period = 0;
    pism_overrides:ocean.delta_mass_flux.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.delta_mass_flux.period_option = "ocean_delta_mass_flux_period";
    pism_overrides:ocean.delta_mass_flux.period_type = "integer";
    pism_overrides:ocean.delta_mass_flux.period_units = "years";

    pism_overrides:ocean.delta_mass_flux.reference_year = 0;
    pism_overrides:ocean.delta_mass_flux.reference_year_doc = "Reference year to use when ``ocean.delta_mass_flux.period`` is active.";
    pism_overrides:ocean.delta_mass_flux.reference_year_option = "ocean_delta_mass_flux_reference_year";
    pism_overrides:ocean.delta_mass_flux.reference_year_type = "integer";
    pism_overrides:ocean.delta_mass_flux.reference_year_units = "years";

    pism_overrides:ocean.delta_sl.file = "";
    pism_overrides:ocean.delta_sl.file_doc = "Name of the file containing sea level offsets.";
    pism_overrides:ocean.delta_sl.file_option = "ocean_delta_sl_file";
    pism_overrides:ocean.delta_sl.file_type = "string";

    pism_overrides:ocean.delta_sl.period = 0;
    pism_overrides:ocean.delta_sl.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.delta_sl.period_option = "ocean_delta_sl_period";
    pism_overrides:ocean.delta_sl.period_type = "integer";
    pism_overrides:ocean.delta_sl.period_units = "years";

    pism_overrides:ocean.delta_sl.reference_year = 0;
    pism_overrides:ocean.delta_sl.reference_year_doc = "Reference year to use when ``ocean.delta_sl.period`` is active.";
    pism_overrides:ocean.delta_sl.reference_year_option = "ocean_delta_sl_reference_year";
    pism_overrides:ocean.delta_sl.reference_year_type = "integer";
    pism_overrides:ocean.delta_sl.reference_year_units = "years";

    pism_overrides:ocean.delta_sl_2d.file = "";
    pism_overrides:ocean.delta_sl_2d.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.delta_sl_2d.file_type = "string";

    pism_overrides:ocean.delta_sl_2d.period = 0;
    pism_overrides:ocean.delta_sl_2d.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.delta_sl_2d.period_type = "integer";
    pism_overrides:ocean.delta_sl_2d.period_units = "years";

    pism_overrides:ocean.delta_sl_2d.reference_year = 0;
    pism_overrides:ocean.delta_sl_2d.reference_year_doc = "Reference year to use when ``ocean.delta_sl_2d.period`` is active.";
    pism_overrides:ocean.delta_sl_2d.reference_year_type = "integer";
    pism_overrides:ocean.delta_sl_2d.reference_year_units = "years";

    pism_overrides:ocean.frac_MBP.file = "";
    pism_overrides:ocean.frac_MBP.file_doc = "Name of the file containing melange back-pressure scaling.";
    pism_overrides:ocean.frac_MBP.file_option = "ocean_frac_MBP_file";
    pism_overrides:ocean.frac_MBP.file_type = "string";

    pism_overrides:ocean.frac_MBP.period = 0;
    pism_overrides:ocean.frac_MBP.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.frac_MBP.period_option = "ocean_frac_MBP_period";
    pism_overrides:ocean.frac_MBP.period_type = "integer";
    pism_overrides:ocean.frac_MBP.period_units = "years";

    pism_overrides:ocean.frac_MBP.reference_year = 0;
    pism_overrides:ocean.frac_MBP.reference_year_doc = "Reference year to use when ``ocean.frac_MBP.period`` is active.";
    pism_overrides:ocean.frac_MBP.reference_year_option = "ocean_frac_MBP_reference_year";
    pism_overrides:ocean.frac_MBP.reference_year_type = "integer";
    pism_overrides:ocean.frac_MBP.reference_year_units = "years";

    pism_overrides:ocean.frac_mass_flux.file = "";
    pism_overrides:ocean.frac_mass_flux.file_doc = "Name of the file containing sub-shelf mass flux scaling.";
    pism_overrides:ocean.frac_mass_flux.file_option = "ocean_frac_mass_flux_file";
    pism_overrides:ocean.frac_mass_flux.file_type = "string";

    pism_overrides:ocean.frac_mass_flux.period = 0;
    pism_overrides:ocean.frac_mass_flux.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.frac_mass_flux.period_option = "ocean_frac_mass_flux_period";
    pism_overrides:ocean.frac_mass_flux.period_type = "integer";
    pism_overrides:ocean.frac_mass_flux.period_units = "years";

    pism_overrides:ocean.frac_mass_flux.reference_year = 0;
    pism_overrides:ocean.frac_mass_flux.reference_year_doc = "Reference year to use when ``ocean.frac_mass_flux.period`` is active.";
    pism_overrides:ocean.frac_mass_flux.reference_year_option = "ocean_frac_mass_flux_reference_year";
    pism_overrides:ocean.frac_mass_flux.reference_year_type = "integer";
    pism_overrides:ocean.frac_mass_flux.reference_year_units = "years";

    pism_overrides:ocean.given.file = "";
    pism_overrides:ocean.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.given.file_option = "ocean_given_file";
    pism_overrides:ocean.given.file_type = "string";

    pism_overrides:ocean.given.period = 0;
    pism_overrides:ocean.given.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.given.period_option = "ocean_given_period";
    pism_overrides:ocean.given.period_type = "integer";
    pism_overrides:ocean.given.period_units = "years";

    pism_overrides:ocean.given.reference_year = 0;
    pism_overrides:ocean.given.reference_year_doc = "Reference year to use when ``ocean.given.period`` is active.";
    pism_overrides:ocean.given.reference_year_option = "ocean_given_reference_year";
    pism_overrides:ocean.given.reference_year_type = "integer";
    pism_overrides:ocean.given.reference_year_units = "years";

    pism_overrides:ocean.ismip6.file = "";
    pism_overrides:ocean.ismip6.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.ismip6.file_option = "ocean_ismip6_file";
    pism_overrides:ocean.ismip6.file_type = "string";

    pism_overrides:ocean.ismip6.period = 0;
    pism_overrides:ocean.ismip6.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.ismip6.period_option = "ocean_ismip6_period";
    pism_overrides:ocean.ismip6.period_type = "integer";
    pism_overrides:ocean.ismip6.period_units = "years";

    pism_overrides:ocean.ismip6.reference_year = 0;
    pism_overrides:ocean.ismip6.reference_year_doc = "Reference year to use when ``ocean.ismip6.period`` is active.";
    pism_overrides:ocean.ismip6.reference_year_option = "ocean_ismip6_reference_year";
    pism_overrides:ocean.ismip6.reference_year_type = "integer";
    pism_overrides:ocean.ismip6.reference_year_units = "years";

    pism_overrides:ocean.ismip6nl.file = "";
    pism_overrides:ocean.ismip6nl.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.ismip6nl.file_option = "ocean_ismip6nl_file";
    pism_overrides:ocean.ismip6nl.file_type = "string";

    pism_overrides:ocean.ismip6nl.period = 0;
    pism_overrides:ocean.ismip6nl.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.ismip6nl.period_option = "ocean_ismip6nl_period";
    pism_overrides:ocean.ismip6nl.period_type = "integer";
    pism_overrides:ocean.ismip6nl.period_units = "years";

    pism_overrides:ocean.ismip6nl.reference_year = 0;
    pism_overrides:ocean.ismip6nl.reference_year_doc = "Reference year to use when ``ocean.ismip6nl.period`` is active.";
    pism_overrides:ocean.ismip6nl.reference_year_option = "ocean_ismip6nl_reference_year";
    pism_overrides:ocean.ismip6nl.reference_year_type = "integer";
    pism_overrides:ocean.ismip6nl.reference_year_units = "years";

    pism_overrides:ocean.melange_back_pressure_fraction = 0.0;
    pism_overrides:ocean.melange_back_pressure_fraction_doc = "default melange back pressure fraction";
    pism_overrides:ocean.melange_back_pressure_fraction_type = "number";
    pism_overrides:ocean.melange_back_pressure_fraction_units = "1";

    pism_overrides:ocean.models = "constant";
    pism_overrides:ocean.models_doc = "Comma-separated list of ocean models and modifiers.";
    pism_overrides:ocean.models_option = "ocean";
    pism_overrides:ocean.models_type = "string";

    pism_overrides:ocean.pico.continental_shelf_depth = -800.0;
    pism_overrides:ocean.pico.continental_shelf_depth_doc = "Determines the edge of the continental shelf to calculate mean ocean properties";
    pism_overrides:ocean.pico.continental_shelf_depth_option = "continental_shelf_depth";
    pism_overrides:ocean.pico.continental_shelf_depth_type = "number";
    pism_overrides:ocean.pico.continental_shelf_depth_units = "meters";

    pism_overrides:ocean.pico.exclude_ice_rises = "yes";
    pism_overrides:ocean.pico.exclude_ice_rises_doc = "Exclude ice rises for box calculation in PICO";
    pism_overrides:ocean.pico.exclude_ice_rises_option = "exclude_icerises";
    pism_overrides:ocean.pico.exclude_ice_rises_type = "flag";

    pism_overrides:ocean.pico.file = "";
    pism_overrides:ocean.pico.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.pico.file_option = "ocean_pico_file";
    pism_overrides:ocean.pico.file_type = "string";

    pism_overrides:ocean.pico.heat_exchange_coefficent = 2e-5;
    pism_overrides:ocean.pico.heat_exchange_coefficent_doc = "Turbulent heat exchange coefficient";
    pism_overrides:ocean.pico.heat_exchange_coefficent_option = "gamma_T";
    pism_overrides:ocean.pico.heat_exchange_coefficent_type = "number";
    pism_overrides:ocean.pico.heat_exchange_coefficent_units = "meters second-1";

    pism_overrides:ocean.pico.maximum_ice_rise_area = 1e5;
    pism_overrides:ocean.pico.maximum_ice_rise_area_doc = "Maximum ice rise area. Patches of grounded ice that are bugger than this are treated as continental ice sheets.";
    pism_overrides:ocean.pico.maximum_ice_rise_area_type = "number";
    pism_overrides:ocean.pico.maximum_ice_rise_area_units = "km2";

    pism_overrides:ocean.pico.number_of_boxes = 5;
    pism_overrides:ocean.pico.number_of_boxes_doc = "Default maximum number of boxes (for the largest ice shelves)";
    pism_overrides:ocean.pico.number_of_boxes_option = "number_of_boxes";
    pism_overrides:ocean.pico.number_of_boxes_type = "integer";
    pism_overrides:ocean.pico.number_of_boxes_units = "pure number";

    pism_overrides:ocean.pico.overturning_coefficent = 1e6;
    pism_overrides:ocean.pico.overturning_coefficent_doc = "Overturning stregth coefficient";
    pism_overrides:ocean.pico.overturning_coefficent_option = "overturning_coeff";
    pism_overrides:ocean.pico.overturning_coefficent_type = "number";
    pism_overrides:ocean.pico.overturning_coefficent_units = "meters6 seconds-1 kg-1";

    pism_overrides:ocean.pico.period = 0;
    pism_overrides:ocean.pico.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.pico.period_option = "ocean_pico_period";
    pism_overrides:ocean.pico.period_type = "integer";
    pism_overrides:ocean.pico.period_units = "years";

    pism_overrides:ocean.pico.reference_year = 0;
    pism_overrides:ocean.pico.reference_year_doc = "Reference year to use when ``ocean.pico.period`` is active.";
    pism_overrides:ocean.pico.reference_year_option = "ocean_pico_reference_year";
    pism_overrides:ocean.pico.reference_year_type = "integer";
    pism_overrides:ocean.pico.reference_year_units = "years";

    pism_overrides:ocean.pik_melt_factor = 5e-3;
    pism_overrides:ocean.pik_melt_factor_doc = "dimensionless tuning parameter in the '-ocean pik' ocean heat flux parameterization; see :cite:`Martinetal2011`";
    pism_overrides:ocean.pik_melt_factor_option = "meltfactor_pik";
    pism_overrides:ocean.pik_melt_factor_type = "number";
    pism_overrides:ocean.pik_melt_factor_units = "1";

    pism_overrides:ocean.sub_shelf_heat_flux_into_ice = 0.5;
    pism_overrides:ocean.sub_shelf_heat_flux_into_ice_doc = "= J meter-2 second-1; naively chosen default value for heat from ocean; see comments in pism::ocean::Constant::shelf_base_mass_flux().";
    pism_overrides:ocean.sub_shelf_heat_flux_into_ice_type = "number";
    pism_overrides:ocean.sub_shelf_heat_flux_into_ice_units = "W meter-2";

    pism_overrides:ocean.th.file = "";
    pism_overrides:ocean.th.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:ocean.th.file_option = "ocean_th_file";
    pism_overrides:ocean.th.file_type = "string";

    pism_overrides:ocean.th.period = 0;
    pism_overrides:ocean.th.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:ocean.th.period_option = "ocean_th_period";
    pism_overrides:ocean.th.period_type = "integer";
    pism_overrides:ocean.th.period_units = "years";

    pism_overrides:ocean.th.reference_year = 0;
    pism_overrides:ocean.th.reference_year_doc = "Reference year to use when ``ocean.th.period`` is active.";
    pism_overrides:ocean.th.reference_year_option = "ocean_th_reference_year";
    pism_overrides:ocean.th.reference_year_type = "integer";
    pism_overrides:ocean.th.reference_year_units = "years";

    pism_overrides:ocean.three_equation_model_clip_salinity = "yes";
    pism_overrides:ocean.three_equation_model_clip_salinity_doc = "Clip shelf base salinity so that it is in the range [4, 40] k/kg. See :cite:`HollandJenkins1999`.";
    pism_overrides:ocean.three_equation_model_clip_salinity_option = "clip_shelf_base_salinity";
    pism_overrides:ocean.three_equation_model_clip_salinity_type = "flag";

    pism_overrides:output.ISMIP6 = "false";
    pism_overrides:output.ISMIP6_doc = "Follow ISMIP6 conventions (units, variable names, \"standard names\") when writing output variables.";
    pism_overrides:output.ISMIP6_type = "flag";

    pism_overrides:output.ISMIP6_extra_variables = "lithk,orog,topg,hfgeoubed,acabf,libmassbfgr,libmassbffl,dlithkdt,velsurf,zvelsurf,velbase,zvelbase,velmean,litemptop,litempbotgr,litempbotfl,strbasemag,licalvf,lifmassbf,sftgif,sftgrf,sftflf";
    pism_overrides:output.ISMIP6_extra_variables_doc = "Comma-separated list of fields reported by models participating in ISMIP6 simulations.";
    pism_overrides:output.ISMIP6_extra_variables_type = "string";

    pism_overrides:output.ISMIP6_ts_variables = "lim,limnsw,iareagr,iareafl,tendacabf,tendlibmassbf,tendlibmassbffl,tendlicalvf,tendlifmassbf";
    pism_overrides:output.ISMIP6_ts_variables_doc = "Comma-separated list of scalar variables (time series) reported by models participating in ISMIP6 simulations.";
    pism_overrides:output.ISMIP6_ts_variables_type = "string";

    pism_overrides:output.backup_interval = 1.0;
    pism_overrides:output.backup_interval_doc = "wall-clock time between automatic backups";
    pism_overrides:output.backup_interval_option = "backup_interval";
    pism_overrides:output.backup_interval_type = "number";
    pism_overrides:output.backup_interval_units = "hours";

    pism_overrides:output.backup_size = "small";
    pism_overrides:output.backup_size_choices = "none,small,medium,big_2d,big";
    pism_overrides:output.backup_size_doc = "The 'size' of a backup file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_overrides:output.backup_size_option = "backup_size";
    pism_overrides:output.backup_size_type = "keyword";

    pism_overrides:output.extra.append = "no";
    pism_overrides:output.extra.append_doc = "Append to an existing output file.";
    pism_overrides:output.extra.append_option = "extra_append";
    pism_overrides:output.extra.append_type = "flag";

    pism_overrides:output.extra.file = "";
    pism_overrides:output.extra.file_doc = "Name of the output file containing spatially-variable diagnostics.";
    pism_overrides:output.extra.file_option = "extra_file";
    pism_overrides:output.extra.file_type = "string";

    pism_overrides:output.extra.split = "no";
    pism_overrides:output.extra.split_doc = "Save spatially-variable diagnostics to separate files (one per time record).";
    pism_overrides:output.extra.split_option = "extra_split";
    pism_overrides:output.extra.split_type = "flag";

    pism_overrides:output.extra.stop_missing = "yes";
    pism_overrides:output.extra.stop_missing_doc = "Stop if requested variable is not available instead of warning.";
    pism_overrides:output.extra.stop_missing_option = "extra_stop_missing";
    pism_overrides:output.extra.stop_missing_type = "flag";

    pism_overrides:output.extra.times = "";
    pism_overrides:output.extra.times_doc = "List or a range of times defining reporting intervals for spatially-variable diagnostics.";
    pism_overrides:output.extra.times_option = "extra_times";
    pism_overrides:output.extra.times_type = "string";

    pism_overrides:output.extra.vars = "";
    pism_overrides:output.extra.vars_doc = "Comma-separated list of spatially-variable diagnostics.";
    pism_overrides:output.extra.vars_option = "extra_vars";
    pism_overrides:output.extra.vars_type = "string";

    pism_overrides:output.file_name = "unnamed.nc";
    pism_overrides:output.file_name_doc = "The file to save final model results to.";
    pism_overrides:output.file_name_option = "o";
    pism_overrides:output.file_name_type = "string";

    pism_overrides:output.fill_value = -2e9;
    pism_overrides:output.fill_value_doc = "_FillValue used when saving diagnostic quantities";
    pism_overrides:output.fill_value_type = "number";
    pism_overrides:output.fill_value_units = "none";

    pism_overrides:output.format = "netcdf3";
    pism_overrides:output.format_choices = "netcdf3,netcdf4_parallel,pnetcdf,pio_pnetcdf,pio_netcdf4p,pio_netcdf4c,pio_netcdf";
    pism_overrides:output.format_doc = "The I/O format used for spatial fields; 'netcdf3' is the default, 'netcd4_parallel' is available if PISM was built with parallel NetCDF-4, and 'pnetcdf' is available if PISM was built with PnetCDF.";
    pism_overrides:output.format_option = "o_format";
    pism_overrides:output.format_type = "keyword";

    pism_overrides:output.ice_free_thickness_standard = 10.0;
    pism_overrides:output.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a grid cell is considered ice-free for purposes of reporting glacierized area, volume, etc.";
    pism_overrides:output.ice_free_thickness_standard_type = "number";
    pism_overrides:output.ice_free_thickness_standard_units = "meters";

    pism_overrides:output.pio.base = 0;
    pism_overrides:output.pio.base_doc = "Rank of the first I/O task";
    pism_overrides:output.pio.base_type = "integer";
    pism_overrides:output.pio.base_units = "count";

    pism_overrides:output.pio.n_writers = 1;
    pism_overrides:output.pio.n_writers_doc = "Number of I/O tasks to use";
    pism_overrides:output.pio.n_writers_type = "integer";
    pism_overrides:output.pio.n_writers_units = "count";

    pism_overrides:output.pio.stride = 1;
    pism_overrides:output.pio.stride_doc = "Offset between I/O tasks";
    pism_overrides:output.pio.stride_type = "integer";
    pism_overrides:output.pio.stride_units = "count";

    pism_overrides:output.runtime.area_scale_factor_log10 = 6;
    pism_overrides:output.runtime.area_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for area (in km^2) in summary line to stdout";
    pism_overrides:output.runtime.area_scale_factor_log10_option = "summary_area_scale_factor_log10";
    pism_overrides:output.runtime.area_scale_factor_log10_type = "integer";
    pism_overrides:output.runtime.area_scale_factor_log10_units = "pure number";

    pism_overrides:output.runtime.time_unit_name = "year";
    pism_overrides:output.runtime.time_unit_name_doc = "Time units used when printing model time, time step, and maximum horizontal velocity at summary to stdout.  Must be valid udunits for time.  (E.g. choose from year,month,day,hour,minute,second.)";
    pism_overrides:output.runtime.time_unit_name_type = "string";

    pism_overrides:output.runtime.time_use_calendar = "yes";
    pism_overrides:output.runtime.time_use_calendar_doc = "Whether to use the current calendar when printing model time in summary to stdout.";
    pism_overrides:output.runtime.time_use_calendar_type = "flag";

    pism_overrides:output.runtime.viewer.size = 320;
    pism_overrides:output.runtime.viewer.size_doc = "default diagnostic viewer size (number of pixels of the longer side)";
    pism_overrides:output.runtime.viewer.size_option = "view_size";
    pism_overrides:output.runtime.viewer.size_type = "integer";
    pism_overrides:output.runtime.viewer.size_units = "count";

    pism_overrides:output.runtime.viewer.variables = "";
    pism_overrides:output.runtime.viewer.variables_doc = "comma-separated list of map-plane diagnostic quantities to view at runtime";
    pism_overrides:output.runtime.viewer.variables_option = "view";
    pism_overrides:output.runtime.viewer.variables_type = "string";

    pism_overrides:output.runtime.volume_scale_factor_log10 = 6;
    pism_overrides:output.runtime.volume_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for volume (in km^3) in summary line to stdout";
    pism_overrides:output.runtime.volume_scale_factor_log10_option = "summary_vol_scale_factor_log10";
    pism_overrides:output.runtime.volume_scale_factor_log10_type = "integer";
    pism_overrides:output.runtime.volume_scale_factor_log10_units = "pure number";

    pism_overrides:output.size = "medium";
    pism_overrides:output.size_choices = "none,small,medium,big_2d,big";
    pism_overrides:output.size_doc = "The 'size' of an output file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_overrides:output.size_option = "o_size";
    pism_overrides:output.size_type = "keyword";

    pism_overrides:output.sizes.big = "cts,liqfrac,temp,temp_pa,uvel,vvel,wvel,wvel_rel";
    pism_overrides:output.sizes.big_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables and variables listed in output.sizes.medium and output.sizes.big_2d) if 'big' output size is selected. Does not include fields written by sub-models.";
    pism_overrides:output.sizes.big_type = "string";

    pism_overrides:output.sizes.big_2d = "age,bfrict,bheatflx,bmelt,bwp,bwprel,dbdt,effbwp,enthalpybase,enthalpysurf,flux_divergence,hardav,hydroinput,lat,litho_temp,lon,nuH,rank,tempbase,tempicethk,tempicethk_basal,temppabase,tempsurf,thk,thksmooth,tillphi,topg,velbar,velbase,wallmelt,wvelbase";
    pism_overrides:output.sizes.big_2d_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables and variables listed in output.sizes.medium) if 'big_2d' output size is selected. Does not include fields written by boundary models.";
    pism_overrides:output.sizes.big_2d_type = "string";

    pism_overrides:output.sizes.medium = "bwat,bwatvel,climatic_mass_balance,diffusivity,enthalpy,flux,flux_mag,ice_surface_temp,liqfrac,mask,schoofs_theta,strain_rates,taub_mag,tauc,taud_mag,temp_pa,tillwat,topgsmooth,usurf,velbar_mag,velbase_mag,velsurf,velsurf_mag,wvelsurf";
    pism_overrides:output.sizes.medium_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables) if 'medium' output size (the default) is selected. Does not include fields written by sub-models.";
    pism_overrides:output.sizes.medium_type = "string";

    pism_overrides:output.snapshot.file = "";
    pism_overrides:output.snapshot.file_doc = "Snapshot (output) file name (or prefix, if saving to individual files).";
    pism_overrides:output.snapshot.file_option = "save_file";
    pism_overrides:output.snapshot.file_type = "string";

    pism_overrides:output.snapshot.size = "small";
    pism_overrides:output.snapshot.size_choices = "none,small,medium,big_2d,big";
    pism_overrides:output.snapshot.size_doc = "The 'size' of a snapshot file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_overrides:output.snapshot.size_option = "save_size";
    pism_overrides:output.snapshot.size_type = "keyword";

    pism_overrides:output.snapshot.split = "no";
    pism_overrides:output.snapshot.split_doc = "Save model state snapshots to separate files (one per time record).";
    pism_overrides:output.snapshot.split_option = "save_split";
    pism_overrides:output.snapshot.split_type = "flag";

    pism_overrides:output.snapshot.times = "";
    pism_overrides:output.snapshot.times_doc = "List or a range of times to save model state snapshots at.";
    pism_overrides:output.snapshot.times_option = "save_times";
    pism_overrides:output.snapshot.times_type = "string";

    pism_overrides:output.timeseries.append = "false";
    pism_overrides:output.timeseries.append_doc = "If true, append to the scalar time series output file.";
    pism_overrides:output.timeseries.append_option = "ts_append";
    pism_overrides:output.timeseries.append_type = "flag";

    pism_overrides:output.timeseries.buffer_size = 10000;
    pism_overrides:output.timeseries.buffer_size_doc = "Number of scalar diagnostic time-series records to hold in memory before writing to disk. (PISM writes this many time-series records to reduce I/O costs.) Send the USR2 signal to flush time-series.";
    pism_overrides:output.timeseries.buffer_size_type = "integer";
    pism_overrides:output.timeseries.buffer_size_units = "count";

    pism_overrides:output.timeseries.filename = "";
    pism_overrides:output.timeseries.filename_doc = "Name of the file to save scalar time series to. Leave empty to disable reporting scalar time-series.";
    pism_overrides:output.timeseries.filename_option = "ts_file";
    pism_overrides:output.timeseries.filename_type = "string";

    pism_overrides:output.timeseries.times = "";
    pism_overrides:output.timeseries.times_doc = "List or range of times defining reporting time intervals.";
    pism_overrides:output.timeseries.times_option = "ts_times";
    pism_overrides:output.timeseries.times_type = "string";

    pism_overrides:output.timeseries.variables = "";
    pism_overrides:output.timeseries.variables_doc = "Requested scalar (time-series) diagnostics. Leave empty to save all available diagnostics.";
    pism_overrides:output.timeseries.variables_option = "ts_vars";
    pism_overrides:output.timeseries.variables_type = "string";

    pism_overrides:output.use_MKS = "false";
    pism_overrides:output.use_MKS_doc = "Use MKS units in output files.";
    pism_overrides:output.use_MKS_type = "flag";

    pism_overrides:regional.no_model_strip = 5.0;
    pism_overrides:regional.no_model_strip_doc = "Default width of the 'no model strip' in regional setups.";
    pism_overrides:regional.no_model_strip_option = "no_model_strip";
    pism_overrides:regional.no_model_strip_type = "number";
    pism_overrides:regional.no_model_strip_units = "km";

    pism_overrides:regional.no_model_yield_stress = 1000.0;
    pism_overrides:regional.no_model_yield_stress_doc = "High yield stress used in the 'no_model_mask' area in the regional mode.";
    pism_overrides:regional.no_model_yield_stress_type = "number";
    pism_overrides:regional.no_model_yield_stress_units = "kPa";

    pism_overrides:regional.zero_gradient = "false";
    pism_overrides:regional.zero_gradient_doc = "Use zero ice thickness and ice surface gradient in the no_model_mask area.";
    pism_overrides:regional.zero_gradient_option = "zero_grad_where_no_model";
    pism_overrides:regional.zero_gradient_type = "flag";

    pism_overrides:run_info.institution = "";
    pism_overrides:run_info.institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";
    pism_overrides:run_info.institution_option = "institution";
    pism_overrides:run_info.institution_type = "string";

    pism_overrides:run_info.title = "";
    pism_overrides:run_info.title_doc = "Free-form string containing a concise description of the current run. This string is written to output files as the 'title' global attribute.";
    pism_overrides:run_info.title_option = "title";
    pism_overrides:run_info.title_type = "string";

    pism_overrides:sea_level.models = "constant";
    pism_overrides:sea_level.models_doc = "Comma-separated list of sea level models and modifiers.";
    pism_overrides:sea_level.models_option = "sea_level";
    pism_overrides:sea_level.models_type = "string";

    pism_overrides:stress_balance.calving_front_stress_bc = "no";
    pism_overrides:stress_balance.calving_front_stress_bc_doc = "Apply CFBC condition as in :cite:`Albrechtetal2011`, :cite:`Winkelmannetal2011`.  May only apply to some stress balances; e.g. SSAFD as of May 2011.  If not set then a strength-extension is used, as in :cite:`BBssasliding`.";
    pism_overrides:stress_balance.calving_front_stress_bc_option = "cfbc";
    pism_overrides:stress_balance.calving_front_stress_bc_type = "flag";

    pism_overrides:stress_balance.ice_free_thickness_standard = 10.0;
    pism_overrides:stress_balance.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a cell is considered ice-free for purposes of computing ice velocity distribution.";
    pism_overrides:stress_balance.ice_free_thickness_standard_type = "number";
    pism_overrides:stress_balance.ice_free_thickness_standard_units = "meters";

    pism_overrides:stress_balance.model = "sia";
    pism_overrides:stress_balance.model_choices = "none,prescribed_sliding,weertman_sliding,sia,ssa,prescribed_sliding+sia,weertman_sliding+sia,ssa+sia";
    pism_overrides:stress_balance.model_doc = "Stress balance model";
    pism_overrides:stress_balance.model_option = "stress_balance";
    pism_overrides:stress_balance.model_type = "keyword";

    pism_overrides:stress_balance.prescribed_sliding.file = "";
    pism_overrides:stress_balance.prescribed_sliding.file_doc = "The name of the file containing prescribed sliding velocity (variable names: `ubar`, `vbar`).";
    pism_overrides:stress_balance.prescribed_sliding.file_type = "string";

    pism_overrides:stress_balance.sia.Glen_exponent = 3.0;
    pism_overrides:stress_balance.sia.Glen_exponent_doc = "Glen exponent in ice flow law for SIA";
    pism_overrides:stress_balance.sia.Glen_exponent_option = "sia_n";
    pism_overrides:stress_balance.sia.Glen_exponent_type = "number";
    pism_overrides:stress_balance.sia.Glen_exponent_units = "pure number";

    pism_overrides:stress_balance.sia.bed_smoother.range = 5.0e3;
    pism_overrides:stress_balance.sia.bed_smoother.range_doc = "half-width of smoothing domain for stressbalance::BedSmoother, in implementing :cite:`Schoofbasaltopg2003` bed roughness parameterization for SIA; set value to zero to turn off mechanism";
    pism_overrides:stress_balance.sia.bed_smoother.range_option = "bed_smoother_range";
    pism_overrides:stress_balance.sia.bed_smoother.range_type = "number";
    pism_overrides:stress_balance.sia.bed_smoother.range_units = "meters";

    pism_overrides:stress_balance.sia.bed_smoother.theta_min = 0.0;
    pism_overrides:stress_balance.sia.bed_smoother.theta_min_doc = "minimum value of `\\theta` in :cite:`Schoofbasaltopg2003` bed roughness parameterization for SIA";
    pism_overrides:stress_balance.sia.bed_smoother.theta_min_type = "number";
    pism_overrides:stress_balance.sia.bed_smoother.theta_min_units = "1";

    pism_overrides:stress_balance.sia.e_age_coupling = "no";
    pism_overrides:stress_balance.sia.e_age_coupling_doc = "Couple the SIA enhancement factor to age as in :cite:`Greve`.";
    pism_overrides:stress_balance.sia.e_age_coupling_option = "e_age_coupling";
    pism_overrides:stress_balance.sia.e_age_coupling_type = "flag";

    pism_overrides:stress_balance.sia.enhancement_factor = 1.0;
    pism_overrides:stress_balance.sia.enhancement_factor_doc = "Flow enhancement factor for SIA";
    pism_overrides:stress_balance.sia.enhancement_factor_option = "sia_e";
    pism_overrides:stress_balance.sia.enhancement_factor_type = "number";
    pism_overrides:stress_balance.sia.enhancement_factor_units = "1";

    pism_overrides:stress_balance.sia.enhancement_factor_interglacial = 1.0;
    pism_overrides:stress_balance.sia.enhancement_factor_interglacial_doc = "Flow enhancement factor for SIA; used for ice accumulated during interglacial periods.";
    pism_overrides:stress_balance.sia.enhancement_factor_interglacial_option = "sia_e_interglacial";
    pism_overrides:stress_balance.sia.enhancement_factor_interglacial_type = "number";
    pism_overrides:stress_balance.sia.enhancement_factor_interglacial_units = "1";

    pism_overrides:stress_balance.sia.flow_law = "gpbld";
    pism_overrides:stress_balance.sia.flow_law_choices = "arr,arrwarm,gk,gpbld,hooke,isothermal_glen,pb";
    pism_overrides:stress_balance.sia.flow_law_doc = "The SIA flow law.";
    pism_overrides:stress_balance.sia.flow_law_option = "sia_flow_law";
    pism_overrides:stress_balance.sia.flow_law_type = "keyword";

    pism_overrides:stress_balance.sia.grain_size_age_coupling = "no";
    pism_overrides:stress_balance.sia.grain_size_age_coupling_doc = "Use age of the ice to compute grain size to use with the Goldsby-Kohlstedt :cite:`GoldsbyKohlstedt` flow law";
    pism_overrides:stress_balance.sia.grain_size_age_coupling_option = "grain_size_age_coupling";
    pism_overrides:stress_balance.sia.grain_size_age_coupling_type = "flag";

    pism_overrides:stress_balance.sia.limit_diffusivity = "no";
    pism_overrides:stress_balance.sia.limit_diffusivity_doc = "Limit SIA diffusivity by `stress_balance.sia.max_diffusivity`.";
    pism_overrides:stress_balance.sia.limit_diffusivity_option = "limit_sia_diffusivity";
    pism_overrides:stress_balance.sia.limit_diffusivity_type = "flag";

    pism_overrides:stress_balance.sia.max_diffusivity = 200.0;
    pism_overrides:stress_balance.sia.max_diffusivity_doc = "Maximum allowed diffusivity of the SIA flow. PISM stops with an error message if the SIA diffusivity exceeds this limit.";
    pism_overrides:stress_balance.sia.max_diffusivity_type = "number";
    pism_overrides:stress_balance.sia.max_diffusivity_units = "m2 s-1";

    pism_overrides:stress_balance.sia.surface_gradient_method = "haseloff";
    pism_overrides:stress_balance.sia.surface_gradient_method_choices = "eta,haseloff,mahaffy";
    pism_overrides:stress_balance.sia.surface_gradient_method_doc = "method used for surface gradient calculation at staggered grid points";
    pism_overrides:stress_balance.sia.surface_gradient_method_option = "gradient";
    pism_overrides:stress_balance.sia.surface_gradient_method_type = "keyword";

    pism_overrides:stress_balance.ssa.Glen_exponent = 3.0;
    pism_overrides:stress_balance.ssa.Glen_exponent_doc = "Glen exponent in ice flow law for SSA";
    pism_overrides:stress_balance.ssa.Glen_exponent_option = "ssa_n";
    pism_overrides:stress_balance.ssa.Glen_exponent_type = "number";
    pism_overrides:stress_balance.ssa.Glen_exponent_units = "pure number";

    pism_overrides:stress_balance.ssa.compute_surface_gradient_inward = "no";
    pism_overrides:stress_balance.ssa.compute_surface_gradient_inward_doc = "If yes then use inward first-order differencing in computing surface gradient in the SSA objects.";
    pism_overrides:stress_balance.ssa.compute_surface_gradient_inward_type = "flag";

    pism_overrides:stress_balance.ssa.dirichlet_bc = "no";
    pism_overrides:stress_balance.ssa.dirichlet_bc_doc = "apply SSA velocity Dirichlet boundary condition";
    pism_overrides:stress_balance.ssa.dirichlet_bc_option = "ssa_dirichlet_bc";
    pism_overrides:stress_balance.ssa.dirichlet_bc_type = "flag";

    pism_overrides:stress_balance.ssa.enhancement_factor = 1.0;
    pism_overrides:stress_balance.ssa.enhancement_factor_doc = "Flow enhancement factor for SSA";
    pism_overrides:stress_balance.ssa.enhancement_factor_option = "ssa_e";
    pism_overrides:stress_balance.ssa.enhancement_factor_type = "number";
    pism_overrides:stress_balance.ssa.enhancement_factor_units = "1";

    pism_overrides:stress_balance.ssa.enhancement_factor_interglacial = 1.0;
    pism_overrides:stress_balance.ssa.enhancement_factor_interglacial_doc = "Flow enhancement factor for SSA; used for ice accumulated during interglacial periods.";
    pism_overrides:stress_balance.ssa.enhancement_factor_interglacial_option = "ssa_e_interglacial";
    pism_overrides:stress_balance.ssa.enhancement_factor_interglacial_type = "number";
    pism_overrides:stress_balance.ssa.enhancement_factor_interglacial_units = "1";

    pism_overrides:stress_balance.ssa.epsilon = 1.0e13;
    pism_overrides:stress_balance.ssa.epsilon_doc = "Initial amount of regularization in computation of product of effective viscosity and thickness (`\\nu H`).  This default value for `\\nu H` comes e.g. from a hardness for the Ross ice shelf (`\\bar B`) = 1.9e8 Pa `s^{1/3}` :cite:`MacAyealetal` and a typical strain rate of 0.001 1/year for the Ross ice shelf, giving `\\nu = (\\bar B) / (2 \\cdot 0.001^{2/3})` = 9.49e+14 Pa s ~ 30 MPa year, the value in :cite:`Ritzetal2001`, but with a tiny thickness `H` of about 1 cm.";
    pism_overrides:stress_balance.ssa.epsilon_option = "ssa_eps";
    pism_overrides:stress_balance.ssa.epsilon_type = "number";
    pism_overrides:stress_balance.ssa.epsilon_units = "Pascal second meter";

    pism_overrides:stress_balance.ssa.fd.brutal_sliding = "false";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_doc = "Enhance sliding speed brutally.";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_option = "brutal_sliding";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_type = "flag";

    pism_overrides:stress_balance.ssa.fd.brutal_sliding_scale = 1.0;
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_scale_doc = "Brutal SSA Sliding Scale";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_scale_option = "brutal_sliding_scale";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_scale_type = "number";
    pism_overrides:stress_balance.ssa.fd.brutal_sliding_scale_units = "1";

    pism_overrides:stress_balance.ssa.fd.lateral_drag.enabled = "false";
    pism_overrides:stress_balance.ssa.fd.lateral_drag.enabled_doc = "set viscosity at ice shelf margin next to ice free bedrock as friction parameterization";
    pism_overrides:stress_balance.ssa.fd.lateral_drag.enabled_type = "flag";

    pism_overrides:stress_balance.ssa.fd.lateral_drag.viscosity = 5.0e15;
    pism_overrides:stress_balance.ssa.fd.lateral_drag.viscosity_doc = "Staggered Viscosity used as side friction parameterization.";
    pism_overrides:stress_balance.ssa.fd.lateral_drag.viscosity_option = "nu_bedrock";
    pism_overrides:stress_balance.ssa.fd.lateral_drag.viscosity_type = "number";
    pism_overrides:stress_balance.ssa.fd.lateral_drag.viscosity_units = "Pascal second";

    pism_overrides:stress_balance.ssa.fd.max_iterations = 300;
    pism_overrides:stress_balance.ssa.fd.max_iterations_doc = "Maximum number of Picard iterations for the ice viscosity computation, in the SSAFD object";
    pism_overrides:stress_balance.ssa.fd.max_iterations_option = "ssafd_picard_maxi";
    pism_overrides:stress_balance.ssa.fd.max_iterations_type = "integer";
    pism_overrides:stress_balance.ssa.fd.max_iterations_units = "count";

    pism_overrides:stress_balance.ssa.fd.max_speed = 300000;
    pism_overrides:stress_balance.ssa.fd.max_speed_doc = "Upper bound for the ice speed computed by the SSAFD solver.";
    pism_overrides:stress_balance.ssa.fd.max_speed_option = "ssafd_max_speed";
    pism_overrides:stress_balance.ssa.fd.max_speed_type = "number";
    pism_overrides:stress_balance.ssa.fd.max_speed_units = "km s-1";

    pism_overrides:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation = 0.8;
    pism_overrides:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_doc = "In event of 'Effective viscosity not converged' failure, use outer iteration rule nuH <- nuH + f (nuH - nuH_old), where f is this parameter.";
    pism_overrides:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_option = "ssafd_nuH_iter_failure_underrelaxation";
    pism_overrides:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_type = "number";
    pism_overrides:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_units = "pure number";

    pism_overrides:stress_balance.ssa.fd.relative_convergence = 1.0e-4;
    pism_overrides:stress_balance.ssa.fd.relative_convergence_doc = "Relative change tolerance for the effective viscosity in the SSAFD object";
    pism_overrides:stress_balance.ssa.fd.relative_convergence_option = "ssafd_picard_rtol";
    pism_overrides:stress_balance.ssa.fd.relative_convergence_type = "number";
    pism_overrides:stress_balance.ssa.fd.relative_convergence_units = "1";

    pism_overrides:stress_balance.ssa.fd.replace_zero_diagonal_entries = "yes";
    pism_overrides:stress_balance.ssa.fd.replace_zero_diagonal_entries_doc = "Replace zero diagonal entries in the SSAFD matrix with basal_resistance.beta_ice_free_bedrock to avoid solver failures.";
    pism_overrides:stress_balance.ssa.fd.replace_zero_diagonal_entries_type = "flag";

    pism_overrides:stress_balance.ssa.flow_law = "gpbld";
    pism_overrides:stress_balance.ssa.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb";
    pism_overrides:stress_balance.ssa.flow_law_doc = "The SSA flow law.";
    pism_overrides:stress_balance.ssa.flow_law_option = "ssa_flow_law";
    pism_overrides:stress_balance.ssa.flow_law_type = "keyword";

    pism_overrides:stress_balance.ssa.method = "fd";
    pism_overrides:stress_balance.ssa.method_choices = "fd,fem";
    pism_overrides:stress_balance.ssa.method_doc = "Algorithm for computing the SSA solution.";
    pism_overrides:stress_balance.ssa.method_option = "ssa_method";
    pism_overrides:stress_balance.ssa.method_type = "keyword";

    pism_overrides:stress_balance.ssa.read_initial_guess = "yes";
    pism_overrides:stress_balance.ssa.read_initial_guess_doc = "Read the initial guess from the input file when re-starting.";
    pism_overrides:stress_balance.ssa.read_initial_guess_option = "ssa_read_initial_guess";
    pism_overrides:stress_balance.ssa.read_initial_guess_type = "flag";

    pism_overrides:stress_balance.ssa.strength_extension.constant_nu = 9.48680701906572e+14;
    pism_overrides:stress_balance.ssa.strength_extension.constant_nu_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  This value for nu comes from hardness (bar B)=1.9e8 `Pa s^{1/3}` :cite:`MacAyealetal` and a typical strain rate of 0.001 year-1:  `\\nu = (\\bar B) / (2 \\cdot 0.001^{2/3})`.  Compare the value of 9.45e14 Pa s = 30 MPa year in :cite:`Ritzetal2001`.";
    pism_overrides:stress_balance.ssa.strength_extension.constant_nu_type = "number";
    pism_overrides:stress_balance.ssa.strength_extension.constant_nu_units = "Pascal second";

    pism_overrides:stress_balance.ssa.strength_extension.min_thickness = 50.0;
    pism_overrides:stress_balance.ssa.strength_extension.min_thickness_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  At ice thicknesses below this value the product nu*H switches from the normal vertical integral to a constant value.  The geometry itself is not affected by this value.";
    pism_overrides:stress_balance.ssa.strength_extension.min_thickness_type = "number";
    pism_overrides:stress_balance.ssa.strength_extension.min_thickness_units = "meters";

    pism_overrides:stress_balance.vertical_velocity_approximation = "centered";
    pism_overrides:stress_balance.vertical_velocity_approximation_choices = "centered,upstream";
    pism_overrides:stress_balance.vertical_velocity_approximation_doc = "Vertical velocity FD approximation. \"Upstream\" uses first-order finite difference to compute u_x and v_y. Uses basal velocity to make decisions.";
    pism_overrides:stress_balance.vertical_velocity_approximation_option = "vertical_velocity_approximation";
    pism_overrides:stress_balance.vertical_velocity_approximation_type = "keyword";

    pism_overrides:stress_balance.weertman_sliding.A = 1.8e-16;
    pism_overrides:stress_balance.weertman_sliding.A_doc = "Sliding parameter in the Weertman-style sliding parameterization :cite:`Tomkin2007`";
    pism_overrides:stress_balance.weertman_sliding.A_type = "number";
    pism_overrides:stress_balance.weertman_sliding.A_units = "Pa-3 year-1 m-2";

    pism_overrides:stress_balance.weertman_sliding.k = 0.2;
    pism_overrides:stress_balance.weertman_sliding.k_doc = "The ratio of the basal water pressure and the ice overburden pressure in the Weertman-style sliding parameterization.";
    pism_overrides:stress_balance.weertman_sliding.k_type = "number";
    pism_overrides:stress_balance.weertman_sliding.k_units = "1";

    pism_overrides:surface.anomaly.file = "";
    pism_overrides:surface.anomaly.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:surface.anomaly.file_option = "surface_anomaly_file";
    pism_overrides:surface.anomaly.file_type = "string";

    pism_overrides:surface.anomaly.period = 0;
    pism_overrides:surface.anomaly.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.anomaly.period_option = "surface_anomaly_period";
    pism_overrides:surface.anomaly.period_type = "integer";
    pism_overrides:surface.anomaly.period_units = "years";

    pism_overrides:surface.anomaly.reference_year = 0;
    pism_overrides:surface.anomaly.reference_year_doc = "Reference year to use when ``surface.anomaly.period`` is active.";
    pism_overrides:surface.anomaly.reference_year_option = "surface_anomaly_reference_year";
    pism_overrides:surface.anomaly.reference_year_type = "integer";
    pism_overrides:surface.anomaly.reference_year_units = "years";

    pism_overrides:surface.cache.update_interval = 10;
    pism_overrides:surface.cache.update_interval_doc = "Update interval (in years) for the `-surface cache` modifier.";
    pism_overrides:surface.cache.update_interval_type = "integer";
    pism_overrides:surface.cache.update_interval_units = "year";

    pism_overrides:surface.delta_T.file = "";
    pism_overrides:surface.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_overrides:surface.delta_T.file_option = "surface_delta_T_file";
    pism_overrides:surface.delta_T.file_type = "string";

    pism_overrides:surface.delta_T.period = 0;
    pism_overrides:surface.delta_T.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.delta_T.period_option = "surface_delta_T_period";
    pism_overrides:surface.delta_T.period_type = "integer";
    pism_overrides:surface.delta_T.period_units = "years";

    pism_overrides:surface.delta_T.reference_year = 0;
    pism_overrides:surface.delta_T.reference_year_doc = "Reference year to use when ``surface.delta_T.period`` is active.";
    pism_overrides:surface.delta_T.reference_year_option = "surface_delta_T_reference_year";
    pism_overrides:surface.delta_T.reference_year_type = "integer";
    pism_overrides:surface.delta_T.reference_year_units = "years";

    pism_overrides:surface.elevation_change.file = "";
    pism_overrides:surface.elevation_change.file_doc = "Name of the file containing the reference surface elevation field (variable ``usurf``).";
    pism_overrides:surface.elevation_change.file_option = "surface_elevation_change_file";
    pism_overrides:surface.elevation_change.file_type = "string";

    pism_overrides:surface.elevation_change.period = 0;
    pism_overrides:surface.elevation_change.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.elevation_change.period_option = "surface_elevation_change_period";
    pism_overrides:surface.elevation_change.period_type = "integer";
    pism_overrides:surface.elevation_change.period_units = "years";

    pism_overrides:surface.elevation_change.reference_year = 0;
    pism_overrides:surface.elevation_change.reference_year_doc = "Reference year to use when ``surface.elevation_change.period`` is active.";
    pism_overrides:surface.elevation_change.reference_year_option = "surface_elevation_change_reference_year";
    pism_overrides:surface.elevation_change.reference_year_type = "integer";
    pism_overrides:surface.elevation_change.reference_year_units = "years";

    pism_overrides:surface.elevation_change.smb.exp_factor = 0;
    pism_overrides:surface.elevation_change.smb.exp_factor_doc = "Exponential for the surface mass balance.";
    pism_overrides:surface.elevation_change.smb.exp_factor_option = "smb_exp_factor";
    pism_overrides:surface.elevation_change.smb.exp_factor_type = "number";
    pism_overrides:surface.elevation_change.smb.exp_factor_units = "Kelvin-1";

    pism_overrides:surface.elevation_change.smb.lapse_rate = 0;
    pism_overrides:surface.elevation_change.smb.lapse_rate_doc = "Lapse rate for the surface mass balance.";
    pism_overrides:surface.elevation_change.smb.lapse_rate_option = "smb_lapse_rate";
    pism_overrides:surface.elevation_change.smb.lapse_rate_type = "number";
    pism_overrides:surface.elevation_change.smb.lapse_rate_units = "(m / year) / km";

    pism_overrides:surface.elevation_change.smb.method = "shift";
    pism_overrides:surface.elevation_change.smb.method_choices = "scale,shift";
    pism_overrides:surface.elevation_change.smb.method_doc = "Choose the SMB adjustment method. ``scale``: use temperature-change-dependent scaling factor. ``shift``: use the SMB lapse rate.";
    pism_overrides:surface.elevation_change.smb.method_option = "smb_adjustment";
    pism_overrides:surface.elevation_change.smb.method_type = "keyword";

    pism_overrides:surface.elevation_change.temperature_lapse_rate = 0;
    pism_overrides:surface.elevation_change.temperature_lapse_rate_doc = "Lapse rate for the temperature at the top of the ice.";
    pism_overrides:surface.elevation_change.temperature_lapse_rate_option = "temp_lapse_rate";
    pism_overrides:surface.elevation_change.temperature_lapse_rate_type = "number";
    pism_overrides:surface.elevation_change.temperature_lapse_rate_units = "K / km";

    pism_overrides:surface.force_to_thickness.alpha = 0.01;
    pism_overrides:surface.force_to_thickness.alpha_doc = "exponential coefficient in force-to-thickness mechanism";
    pism_overrides:surface.force_to_thickness.alpha_option = "force_to_thickness_alpha";
    pism_overrides:surface.force_to_thickness.alpha_type = "number";
    pism_overrides:surface.force_to_thickness.alpha_units = "year-1";

    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor = 1.0;
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_doc = "surface.force_to_thickness.alpha is multiplied by this factor in areas that are ice-free according to the target ice thickness and surface.force_to_thickness.ice_free_thickness_threshold";
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_option = "force_to_thickness_ice_free_alpha_factor";
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_type = "number";
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_units = "1";

    pism_overrides:surface.force_to_thickness.ice_free_thickness_threshold = 1.0;
    pism_overrides:surface.force_to_thickness.ice_free_thickness_threshold_doc = "threshold of ice thickness in the force-to-thickness target field. Used to determine whether to use surface.force_to_thickness.ice_free_alpha_factor.";
    pism_overrides:surface.force_to_thickness.ice_free_thickness_threshold_option = "force_to_thickness_ice_free_thickness_threshold";
    pism_overrides:surface.force_to_thickness.ice_free_thickness_threshold_type = "number";
    pism_overrides:surface.force_to_thickness.ice_free_thickness_threshold_units = "meters";

    pism_overrides:surface.force_to_thickness.start_time = -4.54e9;
    pism_overrides:surface.force_to_thickness.start_time_doc = "Starting time for the \"force to thickness\" modifier; the default is \"start from the creation of the Earth.\"";
    pism_overrides:surface.force_to_thickness.start_time_type = "number";
    pism_overrides:surface.force_to_thickness.start_time_units = "years";

    pism_overrides:surface.force_to_thickness_file = "";
    pism_overrides:surface.force_to_thickness_file_doc = "The name of the file to read the target ice thickness from.";
    pism_overrides:surface.force_to_thickness_file_option = "force_to_thickness_file";
    pism_overrides:surface.force_to_thickness_file_type = "string";

    pism_overrides:surface.given.file = "";
    pism_overrides:surface.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_overrides:surface.given.file_option = "surface_given_file";
    pism_overrides:surface.given.file_type = "string";

    pism_overrides:surface.given.period = 0;
    pism_overrides:surface.given.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.given.period_option = "surface_given_period";
    pism_overrides:surface.given.period_type = "integer";
    pism_overrides:surface.given.period_units = "years";

    pism_overrides:surface.given.reference_year = 0;
    pism_overrides:surface.given.reference_year_doc = "Reference year to use when ``surface.given.period`` is active.";
    pism_overrides:surface.given.reference_year_option = "surface_given_reference_year";
    pism_overrides:surface.given.reference_year_type = "integer";
    pism_overrides:surface.given.reference_year_units = "years";

    pism_overrides:surface.given.smb_max = 91000;
    pism_overrides:surface.given.smb_max_doc = "Maximum climatic mass balance value (used to check input data). Corresponds to 100 m/year ice equivalent.";
    pism_overrides:surface.given.smb_max_type = "number";
    pism_overrides:surface.given.smb_max_units = "kg m-2 year-1";

    pism_overrides:surface.ismip6.file = "";
    pism_overrides:surface.ismip6.file_doc = "Name of the file containing climate forcing anomaly fields.";
    pism_overrides:surface.ismip6.file_option = "surface_ismip6_file";
    pism_overrides:surface.ismip6.file_type = "string";

    pism_overrides:surface.ismip6.period = 0;
    pism_overrides:surface.ismip6.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.ismip6.period_option = "surface_ismip6_period";
    pism_overrides:surface.ismip6.period_type = "integer";
    pism_overrides:surface.ismip6.period_units = "years";

    pism_overrides:surface.ismip6.reference_file = "";
    pism_overrides:surface.ismip6.reference_file_doc = "Name of the file containing reference climate forcing fields.";
    pism_overrides:surface.ismip6.reference_file_option = "surface_ismip6_reference_file";
    pism_overrides:surface.ismip6.reference_file_type = "string";

    pism_overrides:surface.ismip6.reference_year = 0;
    pism_overrides:surface.ismip6.reference_year_doc = "Reference year to use when ``surface.ismip6.period`` is active.";
    pism_overrides:surface.ismip6.reference_year_type = "integer";
    pism_overrides:surface.ismip6.reference_year_units = "years";

    pism_overrides:surface.models = "given";
    pism_overrides:surface.models_doc = "Comma-separated list of surface models and modifiers.";
    pism_overrides:surface.models_option = "surface";
    pism_overrides:surface.models_type = "string";

    pism_overrides:surface.pdd.air_temp_all_precip_as_rain = 275.15;
    pism_overrides:surface.pdd.air_temp_all_precip_as_rain_doc = "threshold temperature above which all precipitation is rain; must exceed surface.pdd.air_temp_all_precip_as_snow to avoid division by zero, because difference is in a denominator";
    pism_overrides:surface.pdd.air_temp_all_precip_as_rain_type = "number";
    pism_overrides:surface.pdd.air_temp_all_precip_as_rain_units = "Kelvin";

    pism_overrides:surface.pdd.air_temp_all_precip_as_snow = 273.15;
    pism_overrides:surface.pdd.air_temp_all_precip_as_snow_doc = "threshold temperature below which all precipitation is snow";
    pism_overrides:surface.pdd.air_temp_all_precip_as_snow_type = "number";
    pism_overrides:surface.pdd.air_temp_all_precip_as_snow_units = "Kelvin";

    pism_overrides:surface.pdd.balance_year_start_day = 94;
    pism_overrides:surface.pdd.balance_year_start_day_doc = "274 day of year for October 1st, beginning of the balance year in northern latitudes.";
    pism_overrides:surface.pdd.balance_year_start_day_type = "integer";
    pism_overrides:surface.pdd.balance_year_start_day_units = "ordinal day number";

    pism_overrides:surface.pdd.factor_ice = 0.00879120879120879;
    pism_overrides:surface.pdd.factor_ice_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`; = (8 mm liquid-water-equivalent) / (pos degree day)";
    pism_overrides:surface.pdd.factor_ice_type = "number";
    pism_overrides:surface.pdd.factor_ice_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.factor_snow = 0.0032967032967033;
    pism_overrides:surface.pdd.factor_snow_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`; = (3 mm liquid-water-equivalent) / (pos degree day)";
    pism_overrides:surface.pdd.factor_snow_type = "number";
    pism_overrides:surface.pdd.factor_snow_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.fausto.T_c = 272.15;
    pism_overrides:surface.pdd.fausto.T_c_doc = "= -1 + 273.15; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.T_c_type = "number";
    pism_overrides:surface.pdd.fausto.T_c_units = "Kelvin";

    pism_overrides:surface.pdd.fausto.T_w = 283.15;
    pism_overrides:surface.pdd.fausto.T_w_doc = "= 10 + 273.15; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.T_w_type = "number";
    pism_overrides:surface.pdd.fausto.T_w_units = "Kelvin";

    pism_overrides:surface.pdd.fausto.beta_ice_c = 0.015;
    pism_overrides:surface.pdd.fausto.beta_ice_c_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.beta_ice_c_type = "number";
    pism_overrides:surface.pdd.fausto.beta_ice_c_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.fausto.beta_ice_w = 0.007;
    pism_overrides:surface.pdd.fausto.beta_ice_w_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.beta_ice_w_type = "number";
    pism_overrides:surface.pdd.fausto.beta_ice_w_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.fausto.beta_snow_c = 0.003;
    pism_overrides:surface.pdd.fausto.beta_snow_c_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.beta_snow_c_type = "number";
    pism_overrides:surface.pdd.fausto.beta_snow_c_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.fausto.beta_snow_w = 0.003;
    pism_overrides:surface.pdd.fausto.beta_snow_w_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.beta_snow_w_type = "number";
    pism_overrides:surface.pdd.fausto.beta_snow_w_units = "meter / (Kelvin day)";

    pism_overrides:surface.pdd.fausto.enabled = "false";
    pism_overrides:surface.pdd.fausto.enabled_doc = "Set PDD parameters using formulas (6) and (7) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.enabled_option = "pdd_fausto";
    pism_overrides:surface.pdd.fausto.enabled_type = "flag";

    pism_overrides:surface.pdd.fausto.latitude_beta_w = 72.0;
    pism_overrides:surface.pdd.fausto.latitude_beta_w_doc = "latitude below which to use warm case, in formula (6) in :cite:`Faustoetal2009`";
    pism_overrides:surface.pdd.fausto.latitude_beta_w_type = "number";
    pism_overrides:surface.pdd.fausto.latitude_beta_w_units = "degree_north";

    pism_overrides:surface.pdd.firn_compaction_to_accumulation_ratio = 0.75;
    pism_overrides:surface.pdd.firn_compaction_to_accumulation_ratio_doc = "How much firn as a fraction of accumulation is turned into ice";
    pism_overrides:surface.pdd.firn_compaction_to_accumulation_ratio_type = "number";
    pism_overrides:surface.pdd.firn_compaction_to_accumulation_ratio_units = "1";

    pism_overrides:surface.pdd.firn_depth_file = "";
    pism_overrides:surface.pdd.firn_depth_file_doc = "The name of the file to read the firn_depth from.";
    pism_overrides:surface.pdd.firn_depth_file_option = "pdd_firn_depth_file";
    pism_overrides:surface.pdd.firn_depth_file_type = "string";

    pism_overrides:surface.pdd.interpret_precip_as_snow = "no";
    pism_overrides:surface.pdd.interpret_precip_as_snow_doc = "Interpret precipitation as snow fall.";
    pism_overrides:surface.pdd.interpret_precip_as_snow_type = "flag";

    pism_overrides:surface.pdd.max_evals_per_year = 52;
    pism_overrides:surface.pdd.max_evals_per_year_doc = "maximum number of times the PDD scheme will ask for air temperature and precipitation to build location-dependent time series for computing (expected) number of positive degree days and snow accumulation; the default means the PDD uses weekly samples of the annual cycle; see also surface.pdd.std_dev";
    pism_overrides:surface.pdd.max_evals_per_year_type = "integer";
    pism_overrides:surface.pdd.max_evals_per_year_units = "count";

    pism_overrides:surface.pdd.method = "expectation_integral";
    pism_overrides:surface.pdd.method_choices = "expectation_integral,repeatable_random_process,random_process";
    pism_overrides:surface.pdd.method_doc = "PDD implementation method";
    pism_overrides:surface.pdd.method_option = "pdd_method";
    pism_overrides:surface.pdd.method_type = "keyword";

    pism_overrides:surface.pdd.positive_threshold_temp = 273.15;
    pism_overrides:surface.pdd.positive_threshold_temp_doc = "temperature used to determine meaning of 'positive' degree day";
    pism_overrides:surface.pdd.positive_threshold_temp_type = "number";
    pism_overrides:surface.pdd.positive_threshold_temp_units = "Kelvin";

    pism_overrides:surface.pdd.refreeze = 0.6;
    pism_overrides:surface.pdd.refreeze_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`";
    pism_overrides:surface.pdd.refreeze_type = "number";
    pism_overrides:surface.pdd.refreeze_units = "1";

    pism_overrides:surface.pdd.refreeze_ice_melt = "yes";
    pism_overrides:surface.pdd.refreeze_ice_melt_doc = "If set to 'yes', refreeze surface.pdd.refreeze fraction of melted ice, otherwise all of the melted ice runs off.";
    pism_overrides:surface.pdd.refreeze_ice_melt_type = "flag";

    pism_overrides:surface.pdd.std_dev = 5.0;
    pism_overrides:surface.pdd.std_dev_doc = "std dev of daily temp variation; = EISMINT-Greenland value :cite:`RitzEISMINT`";
    pism_overrides:surface.pdd.std_dev_type = "number";
    pism_overrides:surface.pdd.std_dev_units = "Kelvin";

    pism_overrides:surface.pdd.std_dev.file = "";
    pism_overrides:surface.pdd.std_dev.file_doc = "The name of the file to read `air_temp_sd` (standard deviation of air temperature) from.";
    pism_overrides:surface.pdd.std_dev.file_option = "pdd_sd_file";
    pism_overrides:surface.pdd.std_dev.file_type = "string";

    pism_overrides:surface.pdd.std_dev.period = 0;
    pism_overrides:surface.pdd.std_dev.period_doc = "Length of the period of the climate forcing data. Set to zero to disable.";
    pism_overrides:surface.pdd.std_dev.period_option = "pdd_sd_period";
    pism_overrides:surface.pdd.std_dev.period_type = "integer";
    pism_overrides:surface.pdd.std_dev.period_units = "years";

    pism_overrides:surface.pdd.std_dev.reference_year = 0;
    pism_overrides:surface.pdd.std_dev.reference_year_doc = "Reference year to use when ``surface.pdd.std_dev.period`` is active.";
    pism_overrides:surface.pdd.std_dev.reference_year_option = "pdd_sd_reference_year";
    pism_overrides:surface.pdd.std_dev.reference_year_type = "integer";
    pism_overrides:surface.pdd.std_dev.reference_year_units = "years";

    pism_overrides:surface.pdd.std_dev_lapse_lat_base = 72.0;
    pism_overrides:surface.pdd.std_dev_lapse_lat_base_doc = "std_dev is a function of latitude, with value surface.pdd.std_dev at this latitude; this value only active if surface.pdd.std_dev_lapse_lat_rate is nonzero";
    pism_overrides:surface.pdd.std_dev_lapse_lat_base_type = "number";
    pism_overrides:surface.pdd.std_dev_lapse_lat_base_units = "degree_north";

    pism_overrides:surface.pdd.std_dev_lapse_lat_rate = 0.0;
    pism_overrides:surface.pdd.std_dev_lapse_lat_rate_doc = "std_dev is a function of latitude, with rate of change with respect to latitude given by this constant";
    pism_overrides:surface.pdd.std_dev_lapse_lat_rate_type = "number";
    pism_overrides:surface.pdd.std_dev_lapse_lat_rate_units = "Kelvin / degree_north";

    pism_overrides:surface.pdd.std_dev_param_a = -0.15;
    pism_overrides:surface.pdd.std_dev_param_a_doc = "Parameter a in Sigma = a*T + b, with T in degrees C. Used only if surface.pdd.std_dev_use_param is set to yes.";
    pism_overrides:surface.pdd.std_dev_param_a_type = "number";
    pism_overrides:surface.pdd.std_dev_param_a_units = "pure number";

    pism_overrides:surface.pdd.std_dev_param_b = 0.66;
    pism_overrides:surface.pdd.std_dev_param_b_doc = "Parameter b in Sigma = a*T + b, with T in degrees C. Used only if surface.pdd.std_dev_use_param is set to yes.";
    pism_overrides:surface.pdd.std_dev_param_b_type = "number";
    pism_overrides:surface.pdd.std_dev_param_b_units = "Kelvin";

    pism_overrides:surface.pdd.std_dev_use_param = "no";
    pism_overrides:surface.pdd.std_dev_use_param_doc = "Parameterize standard deviation as a linear function of air temperature over ice-covered grid cells. The region of application is controlled by geometry.ice_free_thickness_standard.";
    pism_overrides:surface.pdd.std_dev_use_param_type = "flag";

    pism_overrides:surface.pressure = 0.0;
    pism_overrides:surface.pressure_doc = "atmospheric pressure; = pressure at ice surface";
    pism_overrides:surface.pressure_type = "number";
    pism_overrides:surface.pressure_units = "Pascal";

    pism_overrides:time.calendar = "365_day";
    pism_overrides:time.calendar_choices = "standard,gregorian,proleptic_gregorian,noleap,365_day,360_day,julian,none";
    pism_overrides:time.calendar_doc = "The calendar to use.";
    pism_overrides:time.calendar_option = "calendar";
    pism_overrides:time.calendar_type = "keyword";

    pism_overrides:time.dimension_name = "time";
    pism_overrides:time.dimension_name_doc = "The name of the time dimension in PISM output files.";
    pism_overrides:time.dimension_name_type = "string";

    pism_overrides:time.eemian_end = -114500.0;
    pism_overrides:time.eemian_end_doc = "End of the Eemian interglacial period. See :cite:`Greve97Greenland`.";
    pism_overrides:time.eemian_end_type = "number";
    pism_overrides:time.eemian_end_units = "years";

    pism_overrides:time.eemian_start = -132000.0;
    pism_overrides:time.eemian_start_doc = "Start of the Eemian interglacial period. See :cite:`Greve97Greenland`.";
    pism_overrides:time.eemian_start_type = "number";
    pism_overrides:time.eemian_start_units = "years";

    pism_overrides:time.holocene_start = -11000.0;
    pism_overrides:time.holocene_start_doc = "Start of the Holocene interglacial period. See :cite:`Greve97Greenland`.";
    pism_overrides:time.holocene_start_type = "number";
    pism_overrides:time.holocene_start_units = "years";

    pism_overrides:time.reference_date = "1-1-1";
    pism_overrides:time.reference_date_doc = "year-month-day; reference date used for calendar computations and in PISM output files";
    pism_overrides:time.reference_date_type = "string";

    pism_overrides:time.run_length = 1000;
    pism_overrides:time.run_length_doc = "Default run length";
    pism_overrides:time.run_length_type = "number";
    pism_overrides:time.run_length_units = "years";

    pism_overrides:time.start_year = 0;
    pism_overrides:time.start_year_doc = "Start year.";
    pism_overrides:time.start_year_type = "number";
    pism_overrides:time.start_year_units = "years";

    pism_overrides:time_stepping.adaptive_ratio = 0.12;
    pism_overrides:time_stepping.adaptive_ratio_doc = "Adaptive time stepping ratio for the explicit scheme for the mass balance equation; :cite:`BBL`, inequality (25)";
    pism_overrides:time_stepping.adaptive_ratio_option = "adapt_ratio";
    pism_overrides:time_stepping.adaptive_ratio_type = "number";
    pism_overrides:time_stepping.adaptive_ratio_units = "1";

    pism_overrides:time_stepping.count_steps = "no";
    pism_overrides:time_stepping.count_steps_doc = "If yes, IceModel::run() will count the number of time steps it took.  Sometimes useful for performance evaluation.  Counts all steps, regardless of whether processes (mass continuity, energy, velocity, ...) occurred within the step.";
    pism_overrides:time_stepping.count_steps_option = "count_steps";
    pism_overrides:time_stepping.count_steps_type = "flag";

    pism_overrides:time_stepping.hit_extra_times = "yes";
    pism_overrides:time_stepping.hit_extra_times_doc = "Modify the time-stepping mechanism to hit times requested using -extra_times.";
    pism_overrides:time_stepping.hit_extra_times_option = "extra_force_output_times";
    pism_overrides:time_stepping.hit_extra_times_type = "flag";

    pism_overrides:time_stepping.hit_multiples = 0.0;
    pism_overrides:time_stepping.hit_multiples_doc = "Hit every X years, where X is specified using this parameter. Use 0 to disable";
    pism_overrides:time_stepping.hit_multiples_option = "timestep_hit_multiples";
    pism_overrides:time_stepping.hit_multiples_type = "number";
    pism_overrides:time_stepping.hit_multiples_units = "years";

    pism_overrides:time_stepping.hit_save_times = "no";
    pism_overrides:time_stepping.hit_save_times_doc = "Modify the time-stepping mechanism to hit times requested using -save_times.";
    pism_overrides:time_stepping.hit_save_times_option = "save_force_output_times";
    pism_overrides:time_stepping.hit_save_times_type = "flag";

    pism_overrides:time_stepping.hit_ts_times = "no";
    pism_overrides:time_stepping.hit_ts_times_doc = "Modify the time-stepping mechanism to hit times requested using -ts_times.";
    pism_overrides:time_stepping.hit_ts_times_type = "flag";

    pism_overrides:time_stepping.maximum_time_step = 60.0;
    pism_overrides:time_stepping.maximum_time_step_doc = "Maximum allowed time step length";
    pism_overrides:time_stepping.maximum_time_step_option = "max_dt";
    pism_overrides:time_stepping.maximum_time_step_type = "number";
    pism_overrides:time_stepping.maximum_time_step_units = "years";

    pism_overrides:time_stepping.skip.enabled = "no";
    pism_overrides:time_stepping.skip.enabled_doc = "Use the temperature, age, and SSA stress balance computation skipping mechanism.";
    pism_overrides:time_stepping.skip.enabled_option = "skip";
    pism_overrides:time_stepping.skip.enabled_type = "flag";

    pism_overrides:time_stepping.skip.max = 10;
    pism_overrides:time_stepping.skip.max_doc = "Number of mass-balance steps, including SIA diffusivity updates, to perform before a the temperature, age, and SSA stress balance computations are done";
    pism_overrides:time_stepping.skip.max_option = "skip_max";
    pism_overrides:time_stepping.skip.max_type = "integer";
    pism_overrides:time_stepping.skip.max_units = "count";

    pism_overrides:long_name = "PISM configuration flags and parameters.";
    pism_overrides:long_name_doc = "The 'long_name' attribute is required by CF conventions. It is not used by PISM itself.";
}
