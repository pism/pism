netcdf pism_config {
    variables:
    byte pism_config;
    // boolean flags:
    pism_config:do_mass_conserve = "yes";

    pism_config:do_temp = "yes";

    pism_config:do_skip = "no";

    pism_config:do_plastic_till = "no";

    pism_config:do_pseudo_plastic_till = "no";

    pism_config:do_superpose = "no";

    pism_config:thermal_bedrock = "true";

    pism_config:do_bed_deformation = "no";

    pism_config:do_bed_iso = "no";

    pism_config:ocean_kill = "false";

    pism_config:floating_ice_killed = "false";

    pism_config:is_dry_simulation = "no";

    pism_config:use_ssa_velocity = "no";

    pism_config:include_bmr_in_continuity = "yes";
    pism_config:include_bmr_in_continuity_doc = "Include basal melt rate in continuity";

    pism_config:use_constant_nuh_for_ssa = "no";

    pism_config:compute_surf_grad_inward_ssa = "no";

    // parameters:
    pism_config:enhancement_factor = 1.0;
    pism_config:enhancement_factor_doc = "Flow enhancement factor";

    pism_config:constant_grain_size = 1.0e-3;

    pism_config:no_spokes_level = 0.0;
    pism_config:no_spokes_level_doc = "iterations of smoothing of Sigma";

    pism_config:start_year = 0;

    pism_config:run_length_years = 1000;
    pism_config:run_length_years_doc = "Default run length, years";

    pism_config:adaptive_timestepping_ratio = 0.12;

    pism_config:initial_age_of_ice_years = 0.0;

    pism_config:maximum_time_step_years = 60.0;
    pism_config:maximum_time_step_years_doc = "Maximum allowed time step length, years";

    pism_config:epsilon_ssa = 1.0e15;
    pism_config:epsilon_ssa_doc = "initial amount of (denominator) regularization in computation of effective viscosity";

    pism_config:tauc = 1e4;
    pism_config:tauc_doc = "yield stress for basal till (plastic or pseudo-plastic model); 10^4 Pa = 0.1 bar";

    pism_config:max_hmelt = 2.0;
    pism_config:max_hmelt_doc = "maximum thickness of the basal melt water layer";

    pism_config:minimum_temperature_for_sliding = 273.0;
    pism_config:minimum_temperature_for_sliding_doc = "Kelvin. Note less than ice.meltingTemp; if above this value then decide to slide";

    pism_config:skip_max = 10;

    pism_config:till_phi = 30.0;
    pism_config:till_phi_doc = "till friction angle, degrees";

    pism_config:till_pw_fraction = 0.95;
    pism_config:till_pw_fraction_doc = "pure number; pore water pressure is this fraction of overburden";

    pism_config:till_c_0 = 0.0;
    pism_config:till_c_0_doc = "Pa; cohesion of till; note Schoof uses zero but Paterson pp 168--169 gives range 0 -- 40 kPa; but Paterson notes that '... all the pairs c_0 and phi in the table would give a yield stress for Ice Stream B that exceeds the basal shear stress there...'";

    pism_config:mu_sliding = 0.0;

    pism_config:bed_def_interval_years = 10.0;
    pism_config:bed_def_interval_years_doc = "Interval between bed deformation updates, years";

    pism_config:max_iterations_ssa = 300;
    pism_config:max_iterations_ssa_doc = "Maximum number of iterations for the ice viscosity computation";

    pism_config:global_min_allowed_temp = 200.0;
    pism_config:global_min_allowed_temp_doc = "Minimum allowed ice temperature, Kelvin";

    pism_config:max_low_temp_count = 10;
    pism_config:max_low_temp_count_doc = "Maximum number of grid points with ice temperature below global_min_allowed_temp.";

    // for next constants, note (VELOCITY/LENGTH)^2  is very close to 10^-27; compare "\epsilon^2/L^2" which
    // appears in formula (4.1) in C. Schoof 2006 "A variational approach to ice streams" J Fluid Mech 556 pp 227--251
    pism_config:plastic_regularization = 0.01;
    pism_config:pseudo_plastic_q = 0.25;

    pism_config:pseudo_plastic_uthreshold = 100.0;
    pism_config:pseudo_plastic_uthreshold_doc = "Units: m/a";

    pism_config:ssa_relative_convergence = 1.0e-4;

    pism_config:beta_shelves_drag_too = 180000.0;
    pism_config:beta_shelves_drag_too_doc = "Pa s m^{-1}, (1/10000) of value stated in Hulbe&MacAyeal1999 for ice stream E";

    // These constants are not used (so far):
    pism_config:seconds_per_year = 3.15569259747e7;
    pism_config:seconds_per_year_doc = "This value should match the one used by UDUNITS (see src/udunits/pismudunits.dat).";

    pism_config:earth_gravity = 9.81;
    pism_config:earth_gravity_doc = "acceleration due to gravity, m/s^2";

    pism_config:pi = 3.14159265358979;

    pism_config:gas_constant_R = 8.31441;
    pism_config:gas_constant_R_doc = "ideal gas constant, J/(mol K)";
}