netcdf delta_T {
dimensions:
  nv = 2 ;
  time = UNLIMITED ; // (4 currently)
variables:
  double nv(nv) ;
  double time(time) ;
    time:units = "common_year since 1-1-1" ;
    time:axis = "T" ;
    time:bounds = "time_bounds" ;
    time:calendar = "365_day" ;
    time:long_name = "time" ;
  double time_bounds(time, nv) ;
  double delta_T(time) ;
    delta_T:units = "kelvin" ;
    delta_T:long_name = "temperature offsets" ;
data:

 time        = 0,  100, 900, 1000;
 time_bounds = 0, 100, 100, 500, 500, 900, 900, 1000;
 delta_T     = 0, -30, -30, 0;
}
