netcdf pism_config {
    variables:
    byte pism_config;
    // boolean flags:
    pism_config:do_mass_conserve = "yes";
    pism_config:do_mass_conserve_doc = "Solve the mass conservation equation";

    pism_config:do_temp = "yes";
    pism_config:do_temp_doc = "Solve energy conservation and age equations";

    pism_config:do_skip = "no";
    pism_config:do_skip_doc = "Use the temperature, age, and SSA stress balance computation skipping mechanism";

    pism_config:do_plastic_till = "no";
    pism_config:do_plastic_till_doc = "Use Schoof’s plastic till model for ice streams at all grounded points on the ice sheet";

    pism_config:do_pseudo_plastic_till = "no";
    pism_config:do_pseudo_plastic_till_doc = "Use the pseudo-plastic till model.";

    pism_config:do_superpose = "no";
    pism_config:do_superpose_doc = "Combine the velocity ﬁelds from the SIA and SSA models as in [\\ref BB]. Only eﬀective if used with -ssa.";

    pism_config:thermal_bedrock = "yes";
    pism_config:thermal_bedrock_doc = "Use the bedrock thermal model";

    pism_config:do_bed_deformation = "no";
    pism_config:do_bed_deformation_doc = "Use a bed defirmation model";

    pism_config:do_bed_iso = "no";
    pism_config:do_bed_iso_doc = "Compute bed deformations by simple pointwise isostasy.";

    pism_config:ocean_kill = "false";
    pism_config:ocean_kill_doc = "If used with input from a NetCDF initialization ﬁle which has ice-free ocean mask (value MASK_FLOATING_OCEAN0=7), will zero out ice thicknesses in areas that were ice-free ocean at time zero. This is calving at the location of the original calving front.";

    pism_config:floating_ice_killed = "false";
    pism_config:floating_ice_killed_doc = "If ice is (or becomes) ﬂoating then it is set to thickness zero. This is calving at the grounding line.";

    pism_config:is_dry_simulation = "no";
    pism_config:is_dry_simulation_doc = "Dry (oceanless) simulation";

    pism_config:use_ssa_velocity = "no";
    pism_config:use_ssa_velocity_doc = "Use the equations of the shallow shelf approximation [\\ref MacAyeal, \\ref Morland, \\ref SchoofStream, \\ref WeisGreveHutter] for ice shelves and dragging ice shelves (%i.e. ice streams) where so-indicated by the mask";

    pism_config:include_bmr_in_continuity = "yes";
    pism_config:include_bmr_in_continuity_doc = "Include basal melt rate in the continuity equation";

    pism_config:use_constant_nuh_for_ssa = "no";
    pism_config:use_constant_nuh_for_ssa_doc = "Compute velocities in ice shelves and streams with a constant value for the product of viscosity \\f$\\nu\\f$ and thickness \\f$H\\f$, obtained from the shelf extension";

    pism_config:compute_surf_grad_inward_ssa = "no";

    // parameters:
    pism_config:enhancement_factor = 1.0;
    pism_config:enhancement_factor_doc = "Flow enhancement factor";

    pism_config:constant_grain_size = 1.0e-3;
    pism_config:constant_grain_size_doc = "Default constant grains size to use with the Goldsby-Kohlstedt [\\ref GoldsbyKohlstedt] flow law, meters";

    pism_config:no_spokes_level = 0.0;
    pism_config:no_spokes_level_doc = "iterations of smoothing of Sigma";

    pism_config:start_year = 0;
    pism_config:start_year_doc = "Model year at which to start the run.";

    pism_config:run_length_years = 1000;
    pism_config:run_length_years_doc = "Default run length, years";

    pism_config:adaptive_timestepping_ratio = 0.12;
    pism_config:adaptive_timestepping_ratio_doc = "Adaptive time stepping ratio for the explicit scheme for the mass balance equation";

    pism_config:initial_age_of_ice_years = 0.0;
    pism_config:initial_age_of_ice_years_doc = "Initial age of ice, years";

    pism_config:maximum_time_step_years = 60.0;
    pism_config:maximum_time_step_years_doc = "Maximum allowed time step length, years";

    pism_config:epsilon_ssa = 1.0e15;
    pism_config:epsilon_ssa_doc = "initial amount of (denominator) regularization in computation of effective viscosity";

    pism_config:tauc = 1e4;
    pism_config:tauc_doc = "yield stress for basal till (plastic or pseudo-plastic model); 10^4 Pa = 0.1 bar";

    pism_config:max_hmelt = 2.0;
    pism_config:max_hmelt_doc = "maximum thickness of the basal melt water layer, meters";

    pism_config:minimum_temperature_for_sliding = 273.0;
    pism_config:minimum_temperature_for_sliding_doc = "Kelvin. Note less than ice.meltingTemp; if above this value then decide to slide";

    pism_config:skip_max = 10;
    pism_config:skip_max_doc = "Number of mass-balance steps, including SIA diﬀusivity updates, to perform before a the temperature, age, and SSA stress balance computations are done";

    pism_config:till_phi = 30.0;
    pism_config:till_phi_doc = "till friction angle, degrees";

    pism_config:till_pw_fraction = 0.95;
    pism_config:till_pw_fraction_doc = "pure number; pore water pressure is this fraction of overburden";

    pism_config:till_c_0 = 0.0;
    pism_config:till_c_0_doc = "Pa; cohesion of till; note Schoof uses zero but Paterson pp 168--169 gives range 0--40 kPa; but Paterson notes that '... all the pairs c_0 and phi in the table would give a yield stress for Ice Stream B that exceeds the basal shear stress there...'";

    pism_config:mu_sliding = 0.0;
    pism_config:mu_sliding_doc = "The sliding law parameter in SIA regions of the ice. <i>This kind of sliding is not recommended, which is why it is turned oﬀ by default.</i>";

    pism_config:bed_def_interval_years = 10.0;
    pism_config:bed_def_interval_years_doc = "Interval between bed deformation updates, years";

    pism_config:max_iterations_ssa = 300;
    pism_config:max_iterations_ssa_doc = "Maximum number of iterations for the ice viscosity computation";

    pism_config:global_min_allowed_temp = 200.0;
    pism_config:global_min_allowed_temp_doc = "Minimum allowed ice temperature, Kelvin";

    pism_config:max_low_temp_count = 10;
    pism_config:max_low_temp_count_doc = "Maximum number of grid points with ice temperature below global_min_allowed_temp.";

    // for next constants, note (VELOCITY/LENGTH)^2  is very close to 10^-27; compare "\epsilon^2/L^2" which
    // appears in formula (4.1) in C. Schoof 2006 "A variational approach to ice streams" J Fluid Mech 556 pp 227--251
    pism_config:plastic_regularization = 0.01;
    pism_config:plastic_regularization_doc = "Set the value of \\f$\\epsilon\\f$ regularization of plastic till; this is the second \\f$\\epsilon\\f$ in formula (4.1) in [\\ref SchoofStream]";

    pism_config:pseudo_plastic_q = 0.25;
    pism_config:pseudo_plastic_q_doc = "The exponent of the pseudo-plastic basal resistance model";

    pism_config:pseudo_plastic_uthreshold = 100.0;
    pism_config:pseudo_plastic_uthreshold_doc = "Units: m/a";

    pism_config:ssa_relative_convergence = 1.0e-4;
    pism_config:ssa_relative_convergence_doc = "Relative change tolerance for the eﬀective viscosity";

    pism_config:beta_shelves_drag_too = 180000.0;
    pism_config:beta_shelves_drag_too_doc = "Pa s m^{-1}, (1/10000) of value stated in [\\ref HulbeMacAyeal] for ice stream E";

    // The default values for the factors come from EISMINT-Greenland, [\\ref RitzEISMINT] .
    pism_config:pdd_factor_snow = 0.003;
    pism_config:pdd_factor_snow_doc = "m K-1 day-1; EISMINT-Greenland value [\\ref RitzEISMINT] ; = (3 mm ice-equivalent) / (pos degree day)";

    pism_config:pdd_factor_ice = 0.008;
    pism_config:pdd_factor_ice_doc = "m K-1 day-1; EISMINT-Greenland value [\\ref RitzEISMINT] ; = (8 mm ice-equivalent) / (pos degree day)";

    pism_config:pdd_refreeze = 0.6;
    pism_config:pdd_refreeze_doc = "[pure fraction]; EISMINT-Greenland value [\\ref RitzEISMINT] ";

    pism_config:pdd_std_dev = 5.0;
    pism_config:pdd_std_dev_doc = "K; std dev of daily temp variation; EISMINT-Greenland value [\\ref RitzEISMINT] ";

    pism_config:snow_temp_d_ma = 314.98;
    pism_config:snow_temp_d_ma_doc = "K; = 41.83+273.15; base temperature for formula (1) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_gamma_ma = -0.006309;
    pism_config:snow_temp_gamma_ma_doc = "K m-1; = -6.309 / 1km; mean slope lapse rate for formula (1) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_c_ma = -0.7189;
    pism_config:snow_temp_c_ma_doc = "K (degN)-1; latitude-dependence coefficient for formula (1) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_kappa_ma = 0.0672;
    pism_config:snow_temp_kappa_ma_doc = "K (degW)-1; longitude-dependence coefficient for formula (1) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_d_mj = 287.85;
    pism_config:snow_temp_d_mj_doc = "K; = 14.70+273.15; base temperature for formula (2) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_gamma_mj = -0.005426;
    pism_config:snow_temp_gamma_mj_doc = "K m-1; = -5.426 / 1km; mean slope lapse rate for formula (2) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_c_mj = -0.1585;
    pism_config:snow_temp_c_mj_doc = "K (degN)-1; latitude-dependence coefficient for formula (2) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_kappa_mj = 0.0518;
    pism_config:snow_temp_kappa_mj_doc = "K (degW)-1; longitude-dependence coefficient for formula (2) in \\ref Faustoetal2009 ";

    pism_config:snow_temp_july_day = 196;
    pism_config:snow_temp_july_day_doc = "day; = Julian day for July 15; used in corrected formula (4) in \\ref Faustoetal2009 ";

    // These constants are not used (so far):
    pism_config:seconds_per_year = 3.15569259747e7;
    pism_config:seconds_per_year_doc = "This value should match the one used by UDUNITS (see src/udunits/pismudunits.dat).";

    pism_config:earth_gravity = 9.81;
    pism_config:earth_gravity_doc = "acceleration due to gravity, m/s^2";

    pism_config:pi = 3.14159265358979;
    pism_config:pi_doc = "ratio of a circle's circumference to its diameter";

    pism_config:gas_constant_R = 8.31441;
    pism_config:gas_constant_R_doc = "ideal gas constant, J/(mol K)";
}
