netcdf gumparams {
    variables:
    byte pism_overrides;

    pism_overrides:standard_gravity = 9.81;
    pism_overrides:standard_gravity_doc = "m s-2; = g";

    pism_overrides:ice_density = 1000.0;
    pism_overrides:ice_density_doc = "kg m-3; 1% Xanthan gum in water has same density as water";

    pism_overrides:bed_smoother_range = -1.0;
    pism_overrides:bed_smoother_range_doc = "m; negative value de-activates bed smoother";

    pism_overrides:bootstrapping_geothermal_flux_value_no_var = 0.0;
    pism_overrides:bootstrapping_geothermal_flux_value_no_var_doc = "W m-2; no geothermal";

    pism_overrides:preliminary_time_step_duration = 0.01;
    pism_overrides:preliminary_time_step_duration_doc = "s; 1 s is a long time, so this is better for starting up";

    pism_overrides:summary_time_unit_name = "second";
    pism_overrides:summary_time_unit_name_doc = "";

    pism_overrides:summary_time_use_calendar = "no";
    pism_overrides:summary_time_use_calendar_doc = "";

    pism_overrides:summary_vol_scale_factor_log10 = -15;
    pism_overrides:summary_vol_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for volume in summary line to stdout; -15 gives volume in cm^3";

    pism_overrides:summary_area_scale_factor_log10 = -10;
    pism_overrides:summary_area_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for area in summary line to stdout; -10 gives area in cm^2";

    pism_overrides:mask_icefree_thickness_standard = 1e-8;
    pism_overrides:mask_icefree_thickness_standard_doc = "m; only if the fluid is less than this is a cell marked as ice free";

    pism_overrides:mask_is_floating_thickness_standard = 1e-8;
    pism_overrides:mask_is_floating_thickness_standard_doc = "m; should not matter";

    pism_overrides:adaptive_timestepping_ratio = 0.08;
    pism_overrides:adaptive_timestepping_ratio_doc = "; compare default 0.12; needs to be smaller because it is more shear-thinning?";

    pism_overrides:Glen_exponent = 5.9;
    pism_overrides:Glen_exponent_doc = "; = n;  Sayag & Worster (2012) give n = 5.9 +- 0.2";

    pism_overrides:ice_softness = 9.7316e-09;  // vs (e.g.) 4e-25 Pa-3 s-1 for ice
    pism_overrides:ice_softness_doc = "Pa-n s-1; = A_0 = B_0^(-n) = (2 x 11.4 Pa s^(1/n))^(-n);  Sayag & Worster (2012) give B_0/2 = tilde mu = 11.4 +- 0.25 Pa s^(1/n)";
}
