netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:stress_balance.sia.bed_smoother_range = 0.;
    pism_overrides:stress_balance.sia.bed_smoother_range_doc = "m; half-width of smoothing domain for PISMBedSmoother, in implementing [@ref Schoofbasaltopg2003] bed roughness parameterization for SIA; set value to zero to turn off mechanism";

    pism_overrides:summary_vol_scale_factor_log10 = 0;
    pism_overrides:summary_vol_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for volume (in km^3) in summary line to stdout";

    pism_overrides:summary_area_scale_factor_log10 = 0;
    pism_overrides:summary_area_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for area (in km^2) in summary line to stdout";

    pism_overrides:energy.drainage_target_water_fraction = 0.02;
    pism_overrides:energy.drainage_target_water_fraction_doc = "; liquid water fraction (omega) above which drainage occurs, but below which there is no drainage; see [@ref AschwandenBuelerKhroulevBlatter]";

    pism_overrides:energy.temperate_ice_enthalpy_conductivity_ratio = 0.001;
    pism_overrides:energy.temperate_ice_enthalpy_conductivity_ratio_doc = "pure number; K in cold ice is multiplied by this fraction to give K0 in [@ref AschwandenBuelerKhroulevBlatter]";

}
