netcdf pism_config {
    variables:
    byte pism_config;

    pism_config:age.enabled = "no";
    pism_config:age.enabled_doc = "Solve age equation (advection equation for ice age).";
    pism_config:age.enabled_option = "age";
    pism_config:age.enabled_type = "boolean";

    pism_config:age.initial_value = 0.0;
    pism_config:age.initial_value_doc = "Initial age of ice";
    pism_config:age.initial_value_type = "scalar";
    pism_config:age.initial_value_units = "years";

    pism_config:atmosphere.fausto_air_temp.c_ma = -0.7189;
    pism_config:atmosphere.fausto_air_temp.c_ma_doc = "latitude-dependence coefficient for formula (1) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.c_ma_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.c_ma_units = "Kelvin / degree_north";

    pism_config:atmosphere.fausto_air_temp.c_mj = -0.1585;
    pism_config:atmosphere.fausto_air_temp.c_mj_doc = "latitude-dependence coefficient for formula (2) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.c_mj_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.c_mj_units = "Kelvin / degree_north";

    pism_config:atmosphere.fausto_air_temp.d_ma = 314.98;
    pism_config:atmosphere.fausto_air_temp.d_ma_doc = "41.83+273.15; base temperature for formula (1) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.d_ma_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.d_ma_units = "Kelvin";

    pism_config:atmosphere.fausto_air_temp.d_mj = 287.85;
    pism_config:atmosphere.fausto_air_temp.d_mj_doc = "= 14.70+273.15; base temperature for formula (2) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.d_mj_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.d_mj_units = "Kelvin";

    pism_config:atmosphere.fausto_air_temp.gamma_ma = -0.006309;
    pism_config:atmosphere.fausto_air_temp.gamma_ma_doc = "= -6.309 / 1km; mean slope lapse rate for formula (1) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.gamma_ma_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.gamma_ma_units = "Kelvin / meter";

    pism_config:atmosphere.fausto_air_temp.gamma_mj = -0.005426;
    pism_config:atmosphere.fausto_air_temp.gamma_mj_doc = "= -5.426 / 1km; mean slope lapse rate for formula (2) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.gamma_mj_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.gamma_mj_units = "Kelvin / meter";

    pism_config:atmosphere.fausto_air_temp.kappa_ma = 0.0672;
    pism_config:atmosphere.fausto_air_temp.kappa_ma_doc = "longitude-dependence coefficient for formula (1) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.kappa_ma_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.kappa_ma_units = "Kelvin / degree_west";

    pism_config:atmosphere.fausto_air_temp.kappa_mj = 0.0518;
    pism_config:atmosphere.fausto_air_temp.kappa_mj_doc = "longitude-dependence coefficient for formula (2) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.kappa_mj_type = "scalar";
    pism_config:atmosphere.fausto_air_temp.kappa_mj_units = "Kelvin / degree_west";

    pism_config:atmosphere.fausto_air_temp.summer_peak_day = 196;
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_doc = "day of year for July 15; used in corrected formula (4) in [@ref Faustoetal2009] ";
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_type = "integer";
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_units = "ordinal day number";

    pism_config:atmosphere.precip_exponential_factor_for_temperature = 0.07041666667;
    pism_config:atmosphere.precip_exponential_factor_for_temperature_doc = "= 0.169/2.4; in SeaRISE-Greenland formula for paleo-precipitation from present; a 7.3\% change of precipitation rate for every one degC of temperature change [@ref Huybrechts02] ";
    pism_config:atmosphere.precip_exponential_factor_for_temperature_type = "scalar";
    pism_config:atmosphere.precip_exponential_factor_for_temperature_units = "Kelvin-1";

    pism_config:basal_resistance.beta_ice_free_bedrock = 1.8e9;
    pism_config:basal_resistance.beta_ice_free_bedrock_doc = "value is for ice stream E from [@ref HulbeMacAyeal]; thus sliding velocity, but we hope it doesn't matter much; at 100 m/year the linear sliding law gives 57040 Pa basal shear stress";
    pism_config:basal_resistance.beta_ice_free_bedrock_type = "scalar";
    pism_config:basal_resistance.beta_ice_free_bedrock_units = "Pascal second meter-1";

    pism_config:basal_resistance.plastic.regularization = 0.01;
    pism_config:basal_resistance.plastic.regularization_doc = "Set the value of @f$\\epsilon@f$ regularization of plastic till; this is the second @f$\\epsilon@f$ in formula (4.1) in [@ref SchoofStream]";
    pism_config:basal_resistance.plastic.regularization_option = "plastic_reg";
    pism_config:basal_resistance.plastic.regularization_type = "scalar";
    pism_config:basal_resistance.plastic.regularization_units = "meter / year";

    pism_config:basal_resistance.pseudo_plastic.enabled = "no";
    pism_config:basal_resistance.pseudo_plastic.enabled_doc = "Use the pseudo-plastic till model (basal sliding law).";
    pism_config:basal_resistance.pseudo_plastic.enabled_option = "pseudo_plastic";
    pism_config:basal_resistance.pseudo_plastic.enabled_type = "boolean";

    pism_config:basal_resistance.pseudo_plastic.q = 0.25;
    pism_config:basal_resistance.pseudo_plastic.q_doc = "The exponent of the pseudo-plastic basal resistance model";
    pism_config:basal_resistance.pseudo_plastic.q_option = "pseudo_plastic_q";
    pism_config:basal_resistance.pseudo_plastic.q_type = "scalar";
    pism_config:basal_resistance.pseudo_plastic.q_units = "pure number";

    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor = -1.0;
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_doc = "divides pseudo-plastic tauc (yield stress) by given factor; this would increase sliding by given factor in absence of membrane stresses; not used if negative or zero; not used by default";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_option = "sliding_scale_factor_reduces_tauc";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_type = "scalar";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_units = "1";

    pism_config:basal_resistance.pseudo_plastic.u_threshold = 100.0;
    pism_config:basal_resistance.pseudo_plastic.u_threshold_doc = "threshold velocity of the pseudo-plastic sliding law";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_option = "pseudo_plastic_uthreshold";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_type = "scalar";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_units = "meter / year";

    pism_config:basal_yield_stress.add_transportable_water = "no";
    pism_config:basal_yield_stress.add_transportable_water_doc = "If 'yes' then the water amount in the transport system is added to tillwat in determining tauc (in the Mohr-Coulomb relation).  Normally only the water in the till is used.";
    pism_config:basal_yield_stress.add_transportable_water_option = "tauc_add_transportable_water";
    pism_config:basal_yield_stress.add_transportable_water_type = "boolean";

    pism_config:basal_yield_stress.constant.value = 2e5;
    pism_config:basal_yield_stress.constant.value_doc = "fill value for yield stress for basal till (plastic or pseudo-plastic model); note 2 x 10^5 Pa = 2.0 bar is quite strong and little sliding should occur without an explicit tauc choice altering this default";
    pism_config:basal_yield_stress.constant.value_option = "tauc";
    pism_config:basal_yield_stress.constant.value_type = "scalar";
    pism_config:basal_yield_stress.constant.value_units = "Pascal";

    pism_config:basal_yield_stress.ice_free_bedrock = 1e6;
    pism_config:basal_yield_stress.ice_free_bedrock_doc = "the 'high' yield stress value used in grounded ice-free areas.";
    pism_config:basal_yield_stress.ice_free_bedrock_option = "high_tauc";
    pism_config:basal_yield_stress.ice_free_bedrock_type = "scalar";
    pism_config:basal_yield_stress.ice_free_bedrock_units = "Pascal";

    pism_config:basal_yield_stress.model = "mohr_coulomb";
    pism_config:basal_yield_stress.model_choices = "constant,mohr_coulomb";
    pism_config:basal_yield_stress.model_doc = "The basal yield stress model to use when sliding is active.";
    pism_config:basal_yield_stress.model_option = "yield_stress";
    pism_config:basal_yield_stress.model_type = "keyword";

    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion = 0.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_doc = "cohesion of till; = c_0 in most references; note Schoof uses zero but Paterson pp 168--169 gives range 0--40 kPa; but Paterson notes that '... all the pairs c_0 and phi in the table would give a yield stress for Ice Stream B that exceeds the basal shear stress there...'";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_option = "till_cohesion";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_units = "Pascal";

    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient = 0.12;
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_doc = "coefficient of compressiblity of till; value from [@ref Tulaczyketal2000]";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_option = "till_compressibility_coefficient";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden = 0.02;
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_doc = "delta in notes; N_0 = delta P_o where P_o is overburden pressure; N_0 is reference (low) value of effective pressure (i.e. normal stress); N_0 scales with overburden pressure unlike [@ref Tulaczyketal2000]; default value from Greenland and Antarctic model runs";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_option = "till_effective_fraction_overburden";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water = 0.1;
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_doc = "If basal_yield_stress.add_transportable_water = yes then the water amount in the transport system is added to tillwat in determining tauc.  Normally only the water in the till is used.  This factor multiplies the logarithm in that formula.";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_option = "till_log_factor_transportable_water";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_units = "meters";

    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default = 30.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_doc = "fill value for till friction angle";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_option = "plastic_phi";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure = 1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_doc = "reference effective pressure N_0; value from [@ref Tulaczyketal2000]";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_units = "Pascal";

    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio = 0.69;
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_doc = "void ratio at reference effective pressure N_0; value from [@ref Tulaczyketal2000]";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_option = "till_reference_void_ratio";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled = "no";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_doc = "If THE OPTION -topg_to_phi IS SET THEN THIS WILL BE SET TO 'yes', and then MohrCoulombYieldStress will initialize the tillphi field using a piece-wise linear function of depth described by four parameters.";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_type = "boolean";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max = 15.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_doc = "upper value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min = 5.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_doc = "lower value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max = 1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_doc = "the elevation at which the upper value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_units = "meters";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min = -1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_doc = "the elevation at which the lower value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_type = "scalar";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_units = "meters";

    pism_config:basal_yield_stress.slippery_grounding_lines = "no";
    pism_config:basal_yield_stress.slippery_grounding_lines_doc = "If yes, at icy grounded locations with bed elevations below sea level, within one cell of floating ice or ice-free ocean, make tauc as low as possible from the Mohr-Coulomb relation.  Specifically, at such locations replace the normally-computed tauc from the Mohr-Coulomb relation, which uses the effective pressure from the modeled amount of water in the till, by the minimum value of tauc from Mohr-Coulomb, i.e. by using the effective pressure corresponding to the maximum amount of till-stored water.  Does not alter the modeled or reported amount of till water, nor does this mechanism affect water conservation.";
    pism_config:basal_yield_stress.slippery_grounding_lines_option = "tauc_slippery_grounding_lines";
    pism_config:basal_yield_stress.slippery_grounding_lines_type = "boolean";

    pism_config:bed_deformation.lc.elastic_model = "no";
    pism_config:bed_deformation.lc.elastic_model_doc = "Use the elastic part of the Lingle-Clark bed deformation model.";
    pism_config:bed_deformation.lc.elastic_model_option = "bed_def_lc_elastic_model";
    pism_config:bed_deformation.lc.elastic_model_type = "boolean";

    pism_config:bed_deformation.mantle_density = 3300.0;
    pism_config:bed_deformation.mantle_density_doc = "half-space (mantle) density used by the bed deformation model. See [@ref LingleClark, @ref BLKfastearth]";
    pism_config:bed_deformation.mantle_density_type = "scalar";
    pism_config:bed_deformation.mantle_density_units = "kg meter-3";

    pism_config:bed_deformation.lithosphere_flexural_rigidity = 5.0e24;
    pism_config:bed_deformation.lithosphere_flexural_rigidity_doc = "lithosphere flexural rigidity used by the bed deformation model. See [@ref LingleClark, @ref BLKfastearth]";
    pism_config:bed_deformation.lithosphere_flexural_rigidity_type = "scalar";
    pism_config:bed_deformation.lithosphere_flexural_rigidity_units = "Newton meter";

    pism_config:bed_deformation.mantle_viscosity = 1.0e21;
    pism_config:bed_deformation.mantle_viscosity_doc = "half-space (mantle) viscosity used by the bed deformation model. See [@ref LingleClark, @ref BLKfastearth]";
    pism_config:bed_deformation.mantle_viscosity_type = "scalar";
    pism_config:bed_deformation.mantle_viscosity_units = "Pascal second";

    pism_config:bed_deformation.model = "none";
    pism_config:bed_deformation.model_choices = "none,iso,lc";
    pism_config:bed_deformation.model_doc = "Selects a bed deformation model to use. 'iso' is point-wise isostasy, 'lc' is the Lingle-Clark model (see [@ref LingleClark], requires FFTW3).";
    pism_config:bed_deformation.model_option = "bed_def";
    pism_config:bed_deformation.model_type = "keyword";

    pism_config:bed_deformation.update_interval = 10.0;
    pism_config:bed_deformation.update_interval_doc = "Interval between bed deformation updates";
    pism_config:bed_deformation.update_interval_type = "scalar";
    pism_config:bed_deformation.update_interval_units = "years";

    pism_config:bed_deformation.bed_topography_delta_file = "";
    pism_config:bed_deformation.bed_topography_delta_file_option = "topg_delta_file";
    pism_config:bed_deformation.bed_topography_delta_file_doc = "The name of the file to read the topg_delta from. This field is added to the bed topography during initialization.";
    pism_config:bed_deformation.bed_topography_delta_file_type = "string";

    pism_config:bed_deformation.bed_uplift_file = "";
    pism_config:bed_deformation.bed_uplift_file_option = "uplift_file";
    pism_config:bed_deformation.bed_uplift_file_doc = "The name of the file to read the uplift (dbdt) from. Leave empty to read it from an input file or a regridding file.";
    pism_config:bed_deformation.bed_uplift_file_type = "string";

    pism_config:bootstrapping.defaults.bed = 1.0;
    pism_config:bootstrapping.defaults.bed_doc = "bed elevation value to use if topg (bedrock_altitude) variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bed_type = "scalar";
    pism_config:bootstrapping.defaults.bed_units = "meters";

    pism_config:bootstrapping.defaults.bmelt = 0.0;
    pism_config:bootstrapping.defaults.bmelt_doc = "basal melt rate value to use if variable bmelt is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bmelt_type = "scalar";
    pism_config:bootstrapping.defaults.bmelt_units = "meter / second";

    pism_config:bootstrapping.defaults.bwat = 0.0;
    pism_config:bootstrapping.defaults.bwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bwat_type = "scalar";
    pism_config:bootstrapping.defaults.bwat_units = "meters";

    pism_config:bootstrapping.defaults.bwp = 0.0;
    pism_config:bootstrapping.defaults.bwp_doc = "basal water pressure value to use if variable bwp is absent in bootstrapping file; most hydrology models do not use this value because bwp is diagnostic";
    pism_config:bootstrapping.defaults.bwp_type = "scalar";
    pism_config:bootstrapping.defaults.bwp_units = "Pascal";

    pism_config:bootstrapping.defaults.enwat = 0.0;
    pism_config:bootstrapping.defaults.enwat_doc = "effective englacial water thickness value to use if variable enwat is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.enwat_type = "scalar";
    pism_config:bootstrapping.defaults.enwat_units = "meters";

    pism_config:bootstrapping.defaults.geothermal_flux = 0.042;
    pism_config:bootstrapping.defaults.geothermal_flux_doc = "geothermal flux value to use if bheatflx variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.geothermal_flux_type = "scalar";
    pism_config:bootstrapping.defaults.geothermal_flux_units = "Watt meter-2";

    pism_config:bootstrapping.defaults.ice_thickness = 0.0;
    pism_config:bootstrapping.defaults.ice_thickness_doc = "thickness value to use if thk (land_ice_thickness) variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.ice_thickness_type = "scalar";
    pism_config:bootstrapping.defaults.ice_thickness_units = "meters";

    pism_config:bootstrapping.defaults.tillwat = 0.0;
    pism_config:bootstrapping.defaults.tillwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.tillwat_type = "scalar";
    pism_config:bootstrapping.defaults.tillwat_units = "meters";

    pism_config:bootstrapping.defaults.uplift = 0.0;
    pism_config:bootstrapping.defaults.uplift_doc = "uplift value to use if dbdt variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.uplift_type = "scalar";
    pism_config:bootstrapping.defaults.uplift_units = "meter / second";

    pism_config:bootstrapping.temperature_heuristic = "smb";
    pism_config:bootstrapping.temperature_heuristic_choices = "smb,quartic_guess";
    pism_config:bootstrapping.temperature_heuristic_doc = "The heuristic to use to initialize ice temperature during bootstrapping: 'sbm' uses the new method using the surface mass balance, surface temperature, and the geothermal flux, 'quartic_guess' uses the old method using the surface temperature and the geothermal flux.";
    pism_config:bootstrapping.temperature_heuristic_option = "boot_temperature_heuristic";
    pism_config:bootstrapping.temperature_heuristic_type = "keyword";

    pism_config:calving.eigen_calving.K = 0.0;
    pism_config:calving.eigen_calving.K_doc = "Set proportionality constant to determine calving rate from strain rates.  Note references [@ref Levermannetal2012, @ref Martinetal2011] use K in range 10^9 to 3 x 10^11 m a, that is, 3 x 10^16 to 10^19 m s.";
    pism_config:calving.eigen_calving.K_option = "eigen_calving_K";
    pism_config:calving.eigen_calving.K_type = "scalar";
    pism_config:calving.eigen_calving.K_units = "meter second";

    pism_config:calving.float_kill.margin_only = "no";
    pism_config:calving.float_kill.margin_only_doc = "Apply float_kill at ice margin cells only.";
    pism_config:calving.float_kill.margin_only_option = "float_kill_margin_only";
    pism_config:calving.float_kill.margin_only_type = "boolean";

    pism_config:calving.float_kill.calve_near_grounding_line = "yes";
    pism_config:calving.float_kill.calve_near_grounding_line_doc = "Calve floating ice near the grounding line.";
    pism_config:calving.float_kill.calve_near_grounding_line_option = "float_kill_calve_near_grounding_line";
    pism_config:calving.float_kill.calve_near_grounding_line_type = "boolean";

    pism_config:calving.front_retreat.wrap_around = "false";
    pism_config:calving.front_retreat.wrap_around_doc = "If true, wrap around domain boundaries. This may be needed in some regional synthetic geometry setups.";
    pism_config:calving.front_retreat.wrap_around_option = "calving_wrap_around";
    pism_config:calving.front_retreat.wrap_around_type = "boolean";

    pism_config:calving.front_retreat.use_cfl = "false";
    pism_config:calving.front_retreat.use_cfl_doc = "apply CFL criterion for eigen-calving rate front retreat";
    pism_config:calving.front_retreat.use_cfl_option = "calving_cfl";
    pism_config:calving.front_retreat.use_cfl_type = "boolean";

    pism_config:calving.methods = "";
    pism_config:calving.methods_doc = "comma-separated list of calving methods; one or more of 'eigen_calving', 'ocean_kill', 'float_kill', 'thickness_calving'";
    pism_config:calving.methods_option = "calving";
    pism_config:calving.methods_type = "string";

    pism_config:calving.thickness_calving.threshold = 50.0;
    pism_config:calving.thickness_calving.threshold_doc = "When terminal ice thickness of floating ice shelf is less than this threshold, it will be calved off.";
    pism_config:calving.thickness_calving.threshold_option = "thickness_calving_threshold";
    pism_config:calving.thickness_calving.threshold_type = "scalar";
    pism_config:calving.thickness_calving.threshold_units = "meters";

    pism_config:calving.thickness_calving.threshold_file = "";
    pism_config:calving.thickness_calving.threshold_file_doc = "Name of the file containing the spatially-variable thickness calving threshold. ";
    pism_config:calving.thickness_calving.threshold_file_option = "thickness_calving_threshold_file";
    pism_config:calving.thickness_calving.threshold_file_type = "string";

    pism_config:calving.vonmises.sigma_max = 1.0e6;
    pism_config:calving.vonmises.sigma_max_doc = "Set maximum tensile stress.  Note references [@ref Morlighem2016] use 1.0e6 Pa.";
    pism_config:calving.vonmises.sigma_max_option = "vonmises_calving_sigma_max";
    pism_config:calving.vonmises.sigma_max_type = "scalar";
    pism_config:calving.vonmises.sigma_max_units = "Pa";

    pism_config:climate_forcing.buffer_size = 60;
    pism_config:climate_forcing.buffer_size_doc = "number of 2D climate forcing records to keep in memory; = 5 years of monthly records";
    pism_config:climate_forcing.buffer_size_type = "integer";
    pism_config:climate_forcing.buffer_size_units = "count";

    pism_config:climate_forcing.evaluations_per_year = 52;
    pism_config:climate_forcing.evaluations_per_year_doc = "length of the time-series used to compute temporal averages of forcing data (such as mean annual temperature)";
    pism_config:climate_forcing.evaluations_per_year_type = "integer";
    pism_config:climate_forcing.evaluations_per_year_units = "count";

    pism_config:constants.fresh_water.density = 1000.0;
    pism_config:constants.fresh_water.density_doc = "density of fresh water";
    pism_config:constants.fresh_water.density_type = "scalar";
    pism_config:constants.fresh_water.density_units = "kg meter-3";

    pism_config:constants.fresh_water.latent_heat_of_fusion = 3.34e5;
    pism_config:constants.fresh_water.latent_heat_of_fusion_doc = "latent heat of fusion for water [@ref AschwandenBlatter]";
    pism_config:constants.fresh_water.latent_heat_of_fusion_type = "scalar";
    pism_config:constants.fresh_water.latent_heat_of_fusion_units = "Joule / kg";

    pism_config:constants.fresh_water.melting_point_temperature = 273.15;
    pism_config:constants.fresh_water.melting_point_temperature_doc = "melting point of pure water";
    pism_config:constants.fresh_water.melting_point_temperature_type = "scalar";
    pism_config:constants.fresh_water.melting_point_temperature_units = "Kelvin";

    pism_config:constants.fresh_water.specific_heat_capacity = 4170.0;
    pism_config:constants.fresh_water.specific_heat_capacity_doc = "at melting point T_0 [@ref AschwandenBlatter]";
    pism_config:constants.fresh_water.specific_heat_capacity_type = "scalar";
    pism_config:constants.fresh_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.ice.beta_Clausius_Clapeyron = 7.9e-8;
    pism_config:constants.ice.beta_Clausius_Clapeyron_doc = "Clausius-Clapeyron constant relating melting temperature and pressure: beta = dT / dP [@ref Luethi2002]";
    pism_config:constants.ice.beta_Clausius_Clapeyron_type = "scalar";
    pism_config:constants.ice.beta_Clausius_Clapeyron_units = "Kelvin / Pascal";

    pism_config:constants.ice.density = 910.0;
    pism_config:constants.ice.density_doc = "= rho_i; density of ice in ice sheet";
    pism_config:constants.ice.density_type = "scalar";
    pism_config:constants.ice.density_units = "kg meter-3";

    pism_config:constants.ice.grain_size = 1.0;
    pism_config:constants.ice.grain_size_doc = "Default constant ice grain size to use with the Goldsby-Kohlstedt [@ref GoldsbyKohlstedt] flow law";
    pism_config:constants.ice.grain_size_option = "ice_grain_size";
    pism_config:constants.ice.grain_size_type = "scalar";
    pism_config:constants.ice.grain_size_units = "mm";

    pism_config:constants.ice.specific_heat_capacity = 2009.0;
    pism_config:constants.ice.specific_heat_capacity_doc = "specific heat capacity of pure ice at melting point T_0";
    pism_config:constants.ice.specific_heat_capacity_type = "scalar";
    pism_config:constants.ice.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.ice.thermal_conductivity = 2.10;
    pism_config:constants.ice.thermal_conductivity_doc = "= W m-1 K-1; thermal conductivity of pure ice";
    pism_config:constants.ice.thermal_conductivity_type = "scalar";
    pism_config:constants.ice.thermal_conductivity_units = "Joule / (meter Kelvin second)";

    pism_config:constants.ideal_gas_constant = 8.31441;
    pism_config:constants.ideal_gas_constant_doc = "ideal gas constant";
    pism_config:constants.ideal_gas_constant_type = "scalar";
    pism_config:constants.ideal_gas_constant_units = "Joule / (mol Kelvin)";

    pism_config:constants.sea_water.density = 1028.0;
    pism_config:constants.sea_water.density_doc = "density of sea water";
    pism_config:constants.sea_water.density_type = "scalar";
    pism_config:constants.sea_water.density_units = "kg meter-3";

    pism_config:constants.sea_water.specific_heat_capacity = 3985.0;
    pism_config:constants.sea_water.specific_heat_capacity_doc = "at 35 psu, value taken from http://www.kayelaby.npl.co.uk/general_physics/2_7/2_7_9.html";
    pism_config:constants.sea_water.specific_heat_capacity_type = "scalar";
    pism_config:constants.sea_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.standard_gravity = 9.81;
    pism_config:constants.standard_gravity_doc = "acceleration due to gravity on Earth geoid";
    pism_config:constants.standard_gravity_type = "scalar";
    pism_config:constants.standard_gravity_units = "meter second-2";

    pism_config:energy.allow_temperature_above_melting = "no";
    pism_config:energy.allow_temperature_above_melting_doc = "If set to 'yes', allow temperatures above the pressure-malting point in the cold mode temperature code. Used by some verifiaction tests.";
    pism_config:energy.allow_temperature_above_melting_type = "boolean";

    pism_config:energy.basal_melt.use_grounded_cell_fraction  = "true";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_doc = "If geometry.grounded_cell_fraction is set, use the fractional floatation mask to interpolate the basal melt rate at the grounding line between grounded and floating values.";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_option  = "subgl_basal_melt";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_type  = "boolean";

    pism_config:energy.bedrock_thermal_conductivity = 3.0;
    pism_config:energy.bedrock_thermal_conductivity_doc = "= W m-1 K-1; for bedrock used in thermal model [@ref RitzEISMINT]";
    pism_config:energy.bedrock_thermal_conductivity_type = "scalar";
    pism_config:energy.bedrock_thermal_conductivity_units = "Joule / (meter Kelvin second)";

    pism_config:energy.bedrock_thermal_density = 3300.0;
    pism_config:energy.bedrock_thermal_density_doc = "for bedrock used in thermal model";
    pism_config:energy.bedrock_thermal_density_type = "scalar";
    pism_config:energy.bedrock_thermal_density_units = "kg meter-3";

    pism_config:energy.bedrock_thermal_specific_heat_capacity = 1000.0;
    pism_config:energy.bedrock_thermal_specific_heat_capacity_doc = "for bedrock used in thermal model [@ref RitzEISMINT]";
    pism_config:energy.bedrock_thermal_specific_heat_capacity_type = "scalar";
    pism_config:energy.bedrock_thermal_specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:energy.drainage_maximum_rate = 1.58443823077064e-09;
    pism_config:energy.drainage_maximum_rate_doc = "0.05 year-1; maximum rate at which liquid water fraction in temperate ice could possibly drain; see [@ref AschwandenBuelerKhroulevBlatter]";
    pism_config:energy.drainage_maximum_rate_type = "scalar";
    pism_config:energy.drainage_maximum_rate_units = "second-1";

    pism_config:energy.drainage_target_water_fraction = 0.01;
    pism_config:energy.drainage_target_water_fraction_doc = "liquid water fraction (omega) above which drainage occurs, but below which there is no drainage; see [@ref AschwandenBuelerKhroulevBlatter]";
    pism_config:energy.drainage_target_water_fraction_type = "scalar";
    pism_config:energy.drainage_target_water_fraction_units = "1";

    pism_config:energy.enabled = "yes";
    pism_config:energy.enabled_doc = "Solve energy conservation equations.";
    pism_config:energy.enabled_type = "boolean";

    pism_config:energy.enthalpy_cold_bulge_max = 60270.0;
    pism_config:energy.enthalpy_cold_bulge_max_doc = "= (2009 J kg-1 K-1) * (30 K); maximum amount by which advection can reduce the enthalpy of a column of ice below its surface enthalpy value";
    pism_config:energy.enthalpy_cold_bulge_max_type = "scalar";
    pism_config:energy.enthalpy_cold_bulge_max_units = "Joule / kg";

    pism_config:energy.max_low_temperature_count = 10;
    pism_config:energy.max_low_temperature_count_doc = "Maximum number of grid points with ice temperature below energy.minimum_allowed_temperature.";
    pism_config:energy.max_low_temperature_count_option = "max_low_temps";
    pism_config:energy.max_low_temperature_count_type = "integer";
    pism_config:energy.max_low_temperature_count_units = "count";

    pism_config:energy.minimum_allowed_temperature = 200.0;
    pism_config:energy.minimum_allowed_temperature_doc = "Minimum allowed ice temperature";
    pism_config:energy.minimum_allowed_temperature_option = "low_temp";
    pism_config:energy.minimum_allowed_temperature_type = "scalar";
    pism_config:energy.minimum_allowed_temperature_units = "Kelvin";

    pism_config:energy.temperate_ice_enthalpy_conductivity_ratio = 0.1;
    pism_config:energy.temperate_ice_enthalpy_conductivity_ratio_doc = "K in cold ice is multiplied by this fraction to give K0 in [@ref AschwandenBuelerKhroulevBlatter]";
    pism_config:energy.temperate_ice_enthalpy_conductivity_ratio_type = "scalar";
    pism_config:energy.temperate_ice_enthalpy_conductivity_ratio_units = "pure number";

    pism_config:energy.temperature_based = "no";
    pism_config:energy.temperature_based_doc = "Use cold ice (i.e. not polythermal) methods.";
    pism_config:energy.temperature_based_type = "boolean";

    pism_config:energy.temperature_dependent_thermal_conductivity = "no";
    pism_config:energy.temperature_dependent_thermal_conductivity_doc = "If yes, use varkenthSystemCtx class in the energy step. It is base on formula (4.37) in [@ref GreveBlatter2009]. Otherwise use enthSystemCtx, which has temperature-independent thermal conductivity set by constant ice.thermal_conductivity.";
    pism_config:energy.temperature_dependent_thermal_conductivity_option = "vark";
    pism_config:energy.temperature_dependent_thermal_conductivity_type = "boolean";

    pism_config:enthalpy_converter.T_reference = 223.15;
    pism_config:enthalpy_converter.T_reference_doc = "= T_0 in enthalpy formulas in [@ref AschwandenBuelerKhroulevBlatter]";
    pism_config:enthalpy_converter.T_reference_type = "scalar";
    pism_config:enthalpy_converter.T_reference_units = "Kelvin";

    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance = 0.001;
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_doc = "Tolerance within which ice is treated as temperate (cold-ice mode and diagnostics).";
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_type = "scalar";
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_units = "Kelvin";

    pism_config:flow_law.Hooke.A = 4.42165e-9;
    pism_config:flow_law.Hooke.A_doc = "A_Hooke = (1/B_0)^n where n=3 and B_0 = 1.928 a^(1/3) Pa. See [@ref Hooke]";
    pism_config:flow_law.Hooke.A_type = "scalar";
    pism_config:flow_law.Hooke.A_units = "Pascal-3 second-1";

    pism_config:flow_law.Hooke.C = 0.16612;
    pism_config:flow_law.Hooke.C_doc = "See [@ref Hooke]";
    pism_config:flow_law.Hooke.C_type = "scalar";
    pism_config:flow_law.Hooke.C_units = "Kelvin^{flow_law.Hooke.k}";

    pism_config:flow_law.Hooke.Q = 7.88e4;
    pism_config:flow_law.Hooke.Q_doc = "Activation energy, see [@ref Hooke]";
    pism_config:flow_law.Hooke.Q_type = "scalar";
    pism_config:flow_law.Hooke.Q_units = "Joule / mol";

    pism_config:flow_law.Hooke.Tr = 273.39;
    pism_config:flow_law.Hooke.Tr_doc = "See [@ref Hooke]";
    pism_config:flow_law.Hooke.Tr_type = "scalar";
    pism_config:flow_law.Hooke.Tr_units = "Kelvin";

    pism_config:flow_law.Hooke.k = 1.17;
    pism_config:flow_law.Hooke.k_doc = "See [@ref Hooke]";
    pism_config:flow_law.Hooke.k_type = "scalar";
    pism_config:flow_law.Hooke.k_units = "pure number";

    pism_config:flow_law.Paterson_Budd.A_cold = 3.61e-13;
    pism_config:flow_law.Paterson_Budd.A_cold_doc = "Paterson-Budd A_cold, see [@ref PatersonBudd]";
    pism_config:flow_law.Paterson_Budd.A_cold_type = "scalar";
    pism_config:flow_law.Paterson_Budd.A_cold_units = "Pascal-3 / second";

    pism_config:flow_law.Paterson_Budd.A_warm = 1.73e3;
    pism_config:flow_law.Paterson_Budd.A_warm_doc = "Paterson-Budd A_warm, see [@ref PatersonBudd]";
    pism_config:flow_law.Paterson_Budd.A_warm_type = "scalar";
    pism_config:flow_law.Paterson_Budd.A_warm_units = "Pascal-3 / second";

    pism_config:flow_law.Paterson_Budd.Q_cold = 6.0e4;
    pism_config:flow_law.Paterson_Budd.Q_cold_doc = "Paterson-Budd Q_cold, see [@ref PatersonBudd]";
    pism_config:flow_law.Paterson_Budd.Q_cold_type = "scalar";
    pism_config:flow_law.Paterson_Budd.Q_cold_units = "Joule / mol";

    pism_config:flow_law.Paterson_Budd.Q_warm = 13.9e4;
    pism_config:flow_law.Paterson_Budd.Q_warm_doc = "Paterson-Budd Q_warm, see [@ref PatersonBudd]";
    pism_config:flow_law.Paterson_Budd.Q_warm_type = "scalar";
    pism_config:flow_law.Paterson_Budd.Q_warm_units = "Joule / mol";

    pism_config:flow_law.Paterson_Budd.T_critical = 263.15;
    pism_config:flow_law.Paterson_Budd.T_critical_doc = "Paterson-Budd critical temperature, see [@ref PatersonBudd]";
    pism_config:flow_law.Paterson_Budd.T_critical_type = "scalar";
    pism_config:flow_law.Paterson_Budd.T_critical_units = "Kelvin";

    pism_config:flow_law.Schoof_regularizing_length = 1000.0;
    pism_config:flow_law.Schoof_regularizing_length_doc = "Regularizing length (Schoof definition)";
    pism_config:flow_law.Schoof_regularizing_length_type = "scalar";
    pism_config:flow_law.Schoof_regularizing_length_units = "km";

    pism_config:flow_law.Schoof_regularizing_velocity = 1.0;
    pism_config:flow_law.Schoof_regularizing_velocity_doc = "Regularizing velocity (Schoof definition)";
    pism_config:flow_law.Schoof_regularizing_velocity_type = "scalar";
    pism_config:flow_law.Schoof_regularizing_velocity_units = "meter / year";

    pism_config:flow_law.gpbld.water_frac_coeff = 181.25;
    pism_config:flow_law.gpbld.water_frac_coeff_doc = "coefficient in Glen-Paterson-Budd flow law for extra dependence of softness on liquid water fraction (omega) [@ref GreveBlatter2009, @ref LliboutryDuval1985]";
    pism_config:flow_law.gpbld.water_frac_coeff_type = "scalar";
    pism_config:flow_law.gpbld.water_frac_coeff_units = "pure number";

    pism_config:flow_law.gpbld.water_frac_observed_limit = 0.01;
    pism_config:flow_law.gpbld.water_frac_observed_limit_doc = "maximum value of liquid water fraction omega for which softness values are parameterized by [@ref LliboutryDuval1985]; used in Glen-Paterson-Budd-Lliboutry-Duval flow law; compare [@ref AschwandenBuelerKhroulevBlatter]";
    pism_config:flow_law.gpbld.water_frac_observed_limit_type = "scalar";
    pism_config:flow_law.gpbld.water_frac_observed_limit_units = "1";

    pism_config:flow_law.isothermal_Glen.ice_softness = 3.1689e-24;
    pism_config:flow_law.isothermal_Glen.ice_softness_doc = "ice softness used by IsothermalGlenIce [@ref EISMINT96]";
    pism_config:flow_law.isothermal_Glen.ice_softness_type = "scalar";
    pism_config:flow_law.isothermal_Glen.ice_softness_units = "Pascal-3 second-1";

    pism_config:fracture_density.constant_fd = "no";
    pism_config:fracture_density.constant_fd_doc = "FIXME";
    pism_config:fracture_density.constant_fd_option = "constant_fd";
    pism_config:fracture_density.constant_fd_type = "boolean";

    pism_config:fracture_density.constant_healing = "no";
    pism_config:fracture_density.constant_healing_doc = "Constant healing";
    pism_config:fracture_density.constant_healing_option = "constant_healing";
    pism_config:fracture_density.constant_healing_type = "boolean";

    pism_config:fracture_density.enabled = "no";
    pism_config:fracture_density.enabled_doc = "Calculation of fracture density according to stresses and strain rate field.";
    pism_config:fracture_density.enabled_option = "fractures";
    pism_config:fracture_density.enabled_type = "boolean";

    pism_config:fracture_density.fd2d_scheme = "no";
    pism_config:fracture_density.fd2d_scheme_doc = "FIXME";
    pism_config:fracture_density.fd2d_scheme_option = "scheme_fd2d";
    pism_config:fracture_density.fd2d_scheme_type = "boolean";

    pism_config:fracture_density.fracture_weighted_healing = "no";
    pism_config:fracture_density.fracture_weighted_healing_doc = "Fracture weighted healing";
    pism_config:fracture_density.fracture_weighted_healing_option = "fracture_weighted_healing";
    pism_config:fracture_density.fracture_weighted_healing_type = "boolean";

    pism_config:fracture_density.include_grounded_ice = "no";
    pism_config:fracture_density.include_grounded_ice_doc = "model fracture density in grounded areas";
    pism_config:fracture_density.include_grounded_ice_option = "do_frac_on_grounded";
    pism_config:fracture_density.include_grounded_ice_type = "boolean";

    pism_config:fracture_density.lefm = "no";
    pism_config:fracture_density.lefm_doc = "FIXME";
    pism_config:fracture_density.lefm_option = "lefm";
    pism_config:fracture_density.lefm_type = "boolean";

    pism_config:fracture_density.max_shear_stress = "no";
    pism_config:fracture_density.max_shear_stress_doc = "Use the max. shear stress criterion.";
    pism_config:fracture_density.max_shear_stress_option = "max_shear";
    pism_config:fracture_density.max_shear_stress_type = "boolean";

    pism_config:fracture_density.phi0 = 0.0;
    pism_config:fracture_density.phi0_doc = "FIXME";
    pism_config:fracture_density.phi0_option = "phi0";
    pism_config:fracture_density.phi0_type = "scalar";
    pism_config:fracture_density.phi0_units = "1";

    pism_config:fracture_density.softening_lower_limit = 1.0;
    pism_config:fracture_density.softening_lower_limit_doc = "epsilon in equation (6) in Albrecht and Levermann, 'Fracture-induced softening for large-scale ice dynamics'";
    pism_config:fracture_density.softening_lower_limit_option = "fracture_softening";
    pism_config:fracture_density.softening_lower_limit_type = "scalar";
    pism_config:fracture_density.softening_lower_limit_units = "1";

    pism_config:fracture_density.write_fields = "no";
    pism_config:fracture_density.write_fields_doc = "Writing of fracture density related fields to nc-file.";
    pism_config:fracture_density.write_fields_option = "write_fd_fields";
    pism_config:fracture_density.write_fields_type = "boolean";

    pism_config:geometry.grounded_cell_fraction  = "false";
    pism_config:geometry.grounded_cell_fraction_doc = "Linear interpolation scheme ('LI' in Gladstone et al. 2010) expanded to two dimensions is used if switched on in order to evaluate the position of the grounding line on a subgrid scale.";
    pism_config:geometry.grounded_cell_fraction_option = "subgl";
    pism_config:geometry.grounded_cell_fraction_type = "boolean";

    pism_config:geometry.ice_free_thickness_standard = 0.01;
    pism_config:geometry.ice_free_thickness_standard_doc = "If ice is thinner than this standard then the mask is set to MASK_ICE_FREE_BEDROCK or MASK_ICE_FREE_OCEAN.";
    pism_config:geometry.ice_free_thickness_standard_type = "scalar";
    pism_config:geometry.ice_free_thickness_standard_units = "meters";

    pism_config:geometry.part_grid.enabled = "no";
    pism_config:geometry.part_grid.enabled_doc = "apply partially filled grid cell scheme";
    pism_config:geometry.part_grid.enabled_option = "part_grid";
    pism_config:geometry.part_grid.enabled_type = "boolean";

    pism_config:geometry.remove_icebergs = "no";
    pism_config:geometry.remove_icebergs_doc = "identify and kill detached ice-shelf areas";
    pism_config:geometry.remove_icebergs_option = "kill_icebergs";
    pism_config:geometry.remove_icebergs_type = "boolean";

    pism_config:geometry.update.enabled = "yes";
    pism_config:geometry.update.enabled_doc = "Solve the mass conservation equation";
    pism_config:geometry.update.enabled_option = "mass";
    pism_config:geometry.update.enabled_type = "boolean";

    pism_config:geometry.update.use_basal_melt_rate = "yes";
    pism_config:geometry.update.use_basal_melt_rate_doc = "Include basal melt rate in the continuity equation";
    pism_config:geometry.update.use_basal_melt_rate_option = "bmr_in_cont";
    pism_config:geometry.update.use_basal_melt_rate_type = "boolean";

    pism_config:grid.allow_extrapolation = "no";
    pism_config:grid.allow_extrapolation_doc = "Allow extrapolation during regridding.";
    pism_config:grid.allow_extrapolation_option = "allow_extrapolation";
    pism_config:grid.allow_extrapolation_type = "boolean";

    pism_config:grid.Lbz = 0;
    pism_config:grid.Lbz_doc = "Thickness of the thermal bedrock layer.";
    pism_config:grid.Lbz_type = "scalar";
    pism_config:grid.Lbz_units = "meters";

    pism_config:grid.Lx = 1500e3;
    pism_config:grid.Lx_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_config:grid.Lx_type = "scalar";
    pism_config:grid.Lx_units = "meters";

    pism_config:grid.Ly = 1500e3;
    pism_config:grid.Ly_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_config:grid.Ly_type = "scalar";
    pism_config:grid.Ly_units = "meters";

    pism_config:grid.Lz = 4000;
    pism_config:grid.Lz_doc = "Height of the computational domain.";
    pism_config:grid.Lz_type = "scalar";
    pism_config:grid.Lz_units = "meters";

    pism_config:grid.Mbz = 1;
    pism_config:grid.Mbz_doc = "Number of thermal bedrock layers; 1 level corresponds to no bedrock.";
    pism_config:grid.Mbz_type = "integer";
    pism_config:grid.Mbz_units = "count";

    pism_config:grid.Mx = 61;
    pism_config:grid.Mx_doc = "Number of grid points in the x direction.";
    pism_config:grid.Mx_option = "Mx";
    pism_config:grid.Mx_type = "integer";
    pism_config:grid.Mx_units = "count";

    pism_config:grid.My = 61;
    pism_config:grid.My_doc = "Number of grid points in the y direction.";
    pism_config:grid.My_option = "My";
    pism_config:grid.My_type = "integer";
    pism_config:grid.My_units = "count";

    pism_config:grid.Mz = 31;
    pism_config:grid.Mz_doc = "Number of vertical grid levels in the ice.";
    pism_config:grid.Mz_type = "integer";
    pism_config:grid.Mz_units = "count";

    pism_config:grid.correct_cell_areas = "yes";
    pism_config:grid.correct_cell_areas_doc = "Compute corrected cell areas using WGS84 datum (for ice area and volume computations).";
    pism_config:grid.correct_cell_areas_type = "boolean";

    pism_config:grid.ice_vertical_spacing = "quadratic";
    pism_config:grid.ice_vertical_spacing_choices = "quadratic,equal";
    pism_config:grid.ice_vertical_spacing_doc = "vertical spacing in the ice";
    pism_config:grid.ice_vertical_spacing_option = "z_spacing";
    pism_config:grid.ice_vertical_spacing_type = "keyword";

    pism_config:grid.lambda = 4.0;
    pism_config:grid.lambda_doc = "Vertical grid spacing parameter. Roughly equal to the factor by which the grid is coarser at an end away from the ice-bedrock interface.";
    pism_config:grid.lambda_type = "scalar";
    pism_config:grid.lambda_units = "pure number";

    pism_config:grid.max_stencil_width = 2;
    pism_config:grid.max_stencil_width_doc = "Maximum width of the finite-difference stencil used in PISM.";
    pism_config:grid.max_stencil_width_type = "integer";
    pism_config:grid.max_stencil_width_units = "count";

    pism_config:grid.periodicity = "xy";
    pism_config:grid.periodicity_choices = "none,x,y,xy";
    pism_config:grid.periodicity_doc = "horizontal grid periodicity";
    pism_config:grid.periodicity_option = "periodicity";
    pism_config:grid.periodicity_type = "keyword";

    pism_config:hydrology.cavitation_opening_coefficient = 0.5;
    pism_config:hydrology.cavitation_opening_coefficient_doc = "c_1 in notes; coefficient of cavitation opening term in evolution of layer thickness in hydrology::Distributed";
    pism_config:hydrology.cavitation_opening_coefficient_option = "hydrology_cavitation_opening_coefficient";
    pism_config:hydrology.cavitation_opening_coefficient_type = "scalar";
    pism_config:hydrology.cavitation_opening_coefficient_units = "meter-1";

    pism_config:hydrology.const_bmelt = 3.168876461e-10;
    pism_config:hydrology.const_bmelt_doc = "default value is equivalent to 1 cm per year of melt; only used if hydrology.use_const_bmelt = 'yes'";
    pism_config:hydrology.const_bmelt_option = "hydrology_const_bmelt";
    pism_config:hydrology.const_bmelt_type = "scalar";
    pism_config:hydrology.const_bmelt_units = "meter / second";

    pism_config:hydrology.creep_closure_coefficient = 0.04;
    pism_config:hydrology.creep_closure_coefficient_doc = "c_2 in notes; coefficient of creep closure term in evolution of layer thickness in hydrology::Distributed";
    pism_config:hydrology.creep_closure_coefficient_option = "hydrology_creep_closure_coefficient";
    pism_config:hydrology.creep_closure_coefficient_type = "scalar";
    pism_config:hydrology.creep_closure_coefficient_units = "pure number";

    pism_config:hydrology.gradient_power_in_flux = 1.5;
    pism_config:hydrology.gradient_power_in_flux_doc = "= beta in notes; power beta in Darcy's law q = - k W^alpha |grad psi|^{beta-2} grad psi, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.gradient_power_in_flux_option = "hydrology_gradient_power_in_flux";
    pism_config:hydrology.gradient_power_in_flux_type = "scalar";
    pism_config:hydrology.gradient_power_in_flux_units = "pure number";

    pism_config:hydrology.hydraulic_conductivity = 0.001;
    pism_config:hydrology.hydraulic_conductivity_doc = "= k in notes; lateral conductivity, in Darcy's law, for subglacial water layer; units depend on powers alpha = hydrology.thickness_power_in_flux and beta = hydrology_potential_gradient_power_in_flux; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.hydraulic_conductivity_option = "hydrology_hydraulic_conductivity";
    pism_config:hydrology.hydraulic_conductivity_type = "scalar";
    pism_config:hydrology.hydraulic_conductivity_units = "m^{2 beta - alpha} s^{2 beta - 3} kg^{1-beta}";

    pism_config:hydrology.maximum_time_step = 1.0;
    pism_config:hydrology.maximum_time_step_doc = "maximum allowed time step length used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.maximum_time_step_type = "scalar";
    pism_config:hydrology.maximum_time_step_units = "years";

    pism_config:hydrology.model = "null";
    pism_config:hydrology.model_choices = "null,routing,distributed";
    pism_config:hydrology.model_doc = "Basal hydrology sub-model.";
    pism_config:hydrology.model_option = "hydrology";
    pism_config:hydrology.model_type = "keyword";

    pism_config:hydrology.null_diffuse_till_water = "no";
    pism_config:hydrology.null_diffuse_till_water_doc = "Diffuse stored till water laterally. See equation (11) of [@ref BBssasliding]"; 
    pism_config:hydrology.null_diffuse_till_water_type = "boolean";

    pism_config:hydrology.null_diffusion_distance = 2e4;
    pism_config:hydrology.null_diffusion_distance_doc = "diffusion distance for till water thickness; see equation (11) in [@ref BBssasliding]; only active if hydrology.null_diffuse_till_water is set";
    pism_config:hydrology.null_diffusion_distance_type = "scalar";
    pism_config:hydrology.null_diffusion_distance_units = "meters";

    pism_config:hydrology.null_diffusion_time = 1000.0;
    pism_config:hydrology.null_diffusion_time_doc = "diffusion time for till water thickness; see equation (11) in [@ref BBssasliding]; only active if hydrology.null_diffuse_till_water is set";
    pism_config:hydrology.null_diffusion_time_type = "scalar";
    pism_config:hydrology.null_diffusion_time_units = "years";

    pism_config:hydrology.null_strip_width = -1.0;
    pism_config:hydrology.null_strip_width_doc = "if negative then mechanism is inactive; width of strip around computational domain in which water velocity and water amount are set to zero; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.null_strip_width_type = "scalar";
    pism_config:hydrology.null_strip_width_units = "meters";

    pism_config:hydrology.regularizing_porosity = 0.01;
    pism_config:hydrology.regularizing_porosity_doc = "phi_0 in notes; regularizes pressure equation by multiplying time derivative term";
    pism_config:hydrology.regularizing_porosity_option = "hydrology_regularizing_porosity";
    pism_config:hydrology.regularizing_porosity_type = "scalar";
    pism_config:hydrology.regularizing_porosity_units = "pure number";

    pism_config:hydrology.roughness_scale = 0.1;
    pism_config:hydrology.roughness_scale_doc = "W_r in notes; roughness scale determining maximum amount of cavitation opening in hydrology::Distributed";
    pism_config:hydrology.roughness_scale_option = "hydrology_roughness_scale";
    pism_config:hydrology.roughness_scale_type = "scalar";
    pism_config:hydrology.roughness_scale_units = "meters";

    pism_config:hydrology.thickness_power_in_flux = 1.25;
    pism_config:hydrology.thickness_power_in_flux_doc = "= alpha in notes; power alpha in Darcy's law q = - k W^alpha |grad psi|^{beta-2} grad psi, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.thickness_power_in_flux_option = "hydrology_thickness_power_in_flux";
    pism_config:hydrology.thickness_power_in_flux_type = "scalar";
    pism_config:hydrology.thickness_power_in_flux_units = "1";

    pism_config:hydrology.tillwat_decay_rate = 3.16887646154128e-11;
    pism_config:hydrology.tillwat_decay_rate_doc = "default value is equivalent to 1 mm per year; rate at which tillwat is reduced to zero, in absence of other effects like input";
    pism_config:hydrology.tillwat_decay_rate_option = "hydrology_tillwat_decay_rate";
    pism_config:hydrology.tillwat_decay_rate_type = "scalar";
    pism_config:hydrology.tillwat_decay_rate_units = "meter / second";

    pism_config:hydrology.tillwat_max = 2.0;
    pism_config:hydrology.tillwat_max_doc = "maximum effective thickness of the water stored in till";
    pism_config:hydrology.tillwat_max_option = "hydrology_tillwat_max";
    pism_config:hydrology.tillwat_max_type = "scalar";
    pism_config:hydrology.tillwat_max_units = "meters";

    pism_config:hydrology.use_const_bmelt = "no";
    pism_config:hydrology.use_const_bmelt_doc = "if 'yes', subglacial hydrology model sees basal melt rate which is constant and given by hydrology.const_bmelt";
    pism_config:hydrology.use_const_bmelt_option = "hydrology_use_const_bmelt";
    pism_config:hydrology.use_const_bmelt_type = "boolean";

    pism_config:inverse.design.cH1     = 0;
    pism_config:inverse.design.cH1_doc = "weight of derivative part of an H1 norm for inversion design variables";
    pism_config:inverse.design.cH1_option = "inv_design_cH1";
    pism_config:inverse.design.cH1_type = "scalar";
    pism_config:inverse.design.cH1_units = "1";

    pism_config:inverse.design.cL2 = 1;
    pism_config:inverse.design.cL2_doc = "weight of derivative-free part of an H1 norm for inversion design variables";
    pism_config:inverse.design.cL2_option = "inv_design_cL2";
    pism_config:inverse.design.cL2_type = "scalar";
    pism_config:inverse.design.cL2_units = "1";

    pism_config:inverse.design.func = "sobolevH1";
    pism_config:inverse.design.func_choices = "sobolevH1,tv";
    pism_config:inverse.design.func_doc = "functional used for inversion design variables";
    pism_config:inverse.design.func_option = "inv_design_func";
    pism_config:inverse.design.func_type = "keyword";

    pism_config:inverse.design.param = "exp";
    pism_config:inverse.design.param_choices = "ident,trunc,square,exp";
    pism_config:inverse.design.param_doc = "parameterization of design variables used during inversion";
    pism_config:inverse.design.param_option = "inv_design_param";
    pism_config:inverse.design.param_type = "keyword";

    pism_config:inverse.design.param_hardav_eps = 1e4;
    pism_config:inverse.design.param_hardav_eps_doc = "tiny vertically-averaged hardness used as a substitute for 0 in some tauc parameterizations";
    pism_config:inverse.design.param_hardav_eps_type = "scalar";
    pism_config:inverse.design.param_hardav_eps_units = "Pascal second^(1/3)";

    pism_config:inverse.design.param_hardav_scale = 1e8;
    pism_config:inverse.design.param_hardav_scale_doc = "typical size of ice hardness";
    pism_config:inverse.design.param_hardav_scale_type = "scalar";
    pism_config:inverse.design.param_hardav_scale_units = "Pascal second^(1/3)";

    pism_config:inverse.design.param_tauc_eps = 100;
    pism_config:inverse.design.param_tauc_eps_doc = "tiny yield stress used as a substitute for 0 in some tauc parameterizations";
    pism_config:inverse.design.param_tauc_eps_type = "scalar";
    pism_config:inverse.design.param_tauc_eps_units = "Pascal";

    pism_config:inverse.design.param_tauc_scale = 100000;
    pism_config:inverse.design.param_tauc_scale_doc = "typical size of yield stresses";
    pism_config:inverse.design.param_tauc_scale_type = "scalar";
    pism_config:inverse.design.param_tauc_scale_units = "Pascal";

    pism_config:inverse.design.param_trunc_hardav0 = 1e6;
    pism_config:inverse.design.param_trunc_hardav0_doc = "transition point of change to linear behaviour for design variable parameterization type 'trunc'";
    pism_config:inverse.design.param_trunc_hardav0_type = "scalar";
    pism_config:inverse.design.param_trunc_hardav0_units = "Pascal second^(1/3)";

    pism_config:inverse.design.param_trunc_tauc0 = 1000;
    pism_config:inverse.design.param_trunc_tauc0_doc = "transition point of change to linear behaviour for design variable parameterization type 'trunc'";
    pism_config:inverse.design.param_trunc_tauc0_type = "scalar";
    pism_config:inverse.design.param_trunc_tauc0_units = "Pascal";

    pism_config:inverse.log_ratio_scale = 10;
    pism_config:inverse.log_ratio_scale_doc = "Reference scale for log-ratio functionals";
    pism_config:inverse.log_ratio_scale_option = "inv_log_ratio_scale";
    pism_config:inverse.log_ratio_scale_type = "scalar";
    pism_config:inverse.log_ratio_scale_units = "pure number";

    pism_config:inverse.ssa.hardav_max = 1e10;
    pism_config:inverse.ssa.hardav_max_doc = "Maximum allowed value of hardav for inversions with bound constraints";
    pism_config:inverse.ssa.hardav_max_type = "scalar";
    pism_config:inverse.ssa.hardav_max_units = "Pascal second^(1/3)";

    pism_config:inverse.ssa.hardav_min = 0;
    pism_config:inverse.ssa.hardav_min_doc = "Minimum allowed value of hardav for inversions with bound constraints";
    pism_config:inverse.ssa.hardav_min_type = "scalar";
    pism_config:inverse.ssa.hardav_min_units = "Pascal second^(1/3)";

    pism_config:inverse.ssa.length_scale = 50e3;
    pism_config:inverse.ssa.length_scale_doc = "typical length scale for rescaling derivative norms";
    pism_config:inverse.ssa.length_scale_type = "scalar";
    pism_config:inverse.ssa.length_scale_units = "meters";

    pism_config:inverse.ssa.method = "tikhonov_lmvm";
    pism_config:inverse.ssa.method_choices = "sd,nlcg,ign,tikhonov_lmvm,tikhonov_cg,tikhonov_blmvm,tikhonov_lcl,tikhonov_gn";
    pism_config:inverse.ssa.method_doc = "algorithm to use for SSA inversions";
    pism_config:inverse.ssa.method_option = "inv_method";
    pism_config:inverse.ssa.method_type = "keyword";

    pism_config:inverse.ssa.tauc_max = 5e7;
    pism_config:inverse.ssa.tauc_max_doc = "Maximum allowed value of tauc for inversions with bound constraints";
    pism_config:inverse.ssa.tauc_max_type = "scalar";
    pism_config:inverse.ssa.tauc_max_units = "Pascal";

    pism_config:inverse.ssa.tauc_min = 0;
    pism_config:inverse.ssa.tauc_min_doc = "Minimum allowed value of tauc for inversions with bound constraints";
    pism_config:inverse.ssa.tauc_min_type = "scalar";
    pism_config:inverse.ssa.tauc_min_units = "Pascal";

    pism_config:inverse.ssa.tv_exponent = 1.2;
    pism_config:inverse.ssa.tv_exponent_doc = "Lebesgue exponent for pseudo-TV norm";
    pism_config:inverse.ssa.tv_exponent_option = "inv_ssa_tv_exponent";
    pism_config:inverse.ssa.tv_exponent_type = "scalar";
    pism_config:inverse.ssa.tv_exponent_units = "pure number";

    pism_config:inverse.ssa.velocity_eps = 0.1;
    pism_config:inverse.ssa.velocity_eps_doc = "tiny size of ice velocities during inversion";
    pism_config:inverse.ssa.velocity_eps_type = "scalar";
    pism_config:inverse.ssa.velocity_eps_units = "meter / year";

    pism_config:inverse.ssa.velocity_scale = 100;
    pism_config:inverse.ssa.velocity_scale_doc = "typical size of ice velocities expected during inversion";
    pism_config:inverse.ssa.velocity_scale_type = "scalar";
    pism_config:inverse.ssa.velocity_scale_units = "meter / year";

    pism_config:inverse.state_func = "meansquare";
    pism_config:inverse.state_func_choices = "meansquare,log_ratio,log_relative";
    pism_config:inverse.state_func_doc = "functional used for inversion design variables";
    pism_config:inverse.state_func_option = "inv_state_func";
    pism_config:inverse.state_func_type = "keyword";

    pism_config:inverse.target_misfit = 100;
    pism_config:inverse.target_misfit_doc = "desired root misfit for SSA inversions";
    pism_config:inverse.target_misfit_option = "inv_target_misfit";
    pism_config:inverse.target_misfit_type = "scalar";
    pism_config:inverse.target_misfit_units = "meter / year";

    pism_config:inverse.tikhonov.atol = 1e-10;
    pism_config:inverse.tikhonov.atol_doc = "absolute threshold for Tikhonov stopping criterion";
    pism_config:inverse.tikhonov.atol_option = "tikhonov_atol";
    pism_config:inverse.tikhonov.atol_type = "scalar";
    pism_config:inverse.tikhonov.atol_units = "meter / year";

    pism_config:inverse.tikhonov.penalty_weight = 1;
    pism_config:inverse.tikhonov.penalty_weight_doc = "penalty parameter for Tikhonov inversion";
    pism_config:inverse.tikhonov.penalty_weight_option = "tikhonov_penalty";
    pism_config:inverse.tikhonov.penalty_weight_type = "scalar";
    pism_config:inverse.tikhonov.penalty_weight_units = "1";

    pism_config:inverse.tikhonov.ptol = 0.1;
    pism_config:inverse.tikhonov.ptol_doc = "threshold for reaching desired misfit for adaptive Tikhonov algorithms";
    pism_config:inverse.tikhonov.ptol_option = "tikhonov_ptol";
    pism_config:inverse.tikhonov.ptol_type = "scalar";
    pism_config:inverse.tikhonov.ptol_units = "pure number";

    pism_config:inverse.tikhonov.rtol = 5e-2;
    pism_config:inverse.tikhonov.rtol_doc = "relative threshold for Tikhonov stopping criterion";
    pism_config:inverse.tikhonov.rtol_option = "tikhonov_rtol";
    pism_config:inverse.tikhonov.rtol_type = "scalar";
    pism_config:inverse.tikhonov.rtol_units = "1";

    pism_config:ocean.always_grounded = "no";
    pism_config:ocean.always_grounded_doc = "Dry (ocean-less) simulation; ice is considered grounded regardless of ice thickness, bed elevation, and sea level.";
    pism_config:ocean.always_grounded_option = "dry";
    pism_config:ocean.always_grounded_type = "boolean";

    pism_config:ocean.pik_melt_factor = 5e-3;
    pism_config:ocean.pik_melt_factor_doc = "dimensionless tuning parameter in the '-ocean pik' ocean heat flux parameterization; see [@ref Martinetal2011]";
    pism_config:ocean.pik_melt_factor_option = "meltfactor_pik";
    pism_config:ocean.pik_melt_factor_type = "scalar";
    pism_config:ocean.pik_melt_factor_units = "1";

    pism_config:ocean.runoff_to_ocean_melt_b = 0.15;
    pism_config:ocean.runoff_to_ocean_melt_b_doc = "parameter B in eqn. 1 in @ref Aschwanden";
    pism_config:ocean.runoff_to_ocean_melt_b_type = "scalar";
    pism_config:ocean.runoff_to_ocean_melt_b_units = "1";

    pism_config:ocean.runoff_to_ocean_melt_power_alpha = 0.54;
    pism_config:ocean.runoff_to_ocean_melt_power_alpha_doc = "exponent alpha in eqn. 1 in @ref Xu2013";
    pism_config:ocean.runoff_to_ocean_melt_power_alpha_type = "scalar";
    pism_config:ocean.runoff_to_ocean_melt_power_alpha_units = "1";

    pism_config:ocean.runoff_to_ocean_melt_power_beta = 1.17;
    pism_config:ocean.runoff_to_ocean_melt_power_beta_doc = "exponent beta in eqn. 1 in @ref Xu2013";
    pism_config:ocean.runoff_to_ocean_melt_power_beta_type = "scalar";
    pism_config:ocean.runoff_to_ocean_melt_power_beta_units = "1";

    pism_config:ocean.sub_shelf_heat_flux_into_ice = 0.5;
    pism_config:ocean.sub_shelf_heat_flux_into_ice_doc = "= J meter-2 second-1; naively chosen default value for heat from ocean; see comments in @ref pism::ocean::Constant::shelf_base_mass_flux().";
    pism_config:ocean.sub_shelf_heat_flux_into_ice_type = "scalar";
    pism_config:ocean.sub_shelf_heat_flux_into_ice_units = "W meter-2";

    pism_config:ocean.three_equation_model_clip_salinity = "yes";
    pism_config:ocean.three_equation_model_clip_salinity_doc = "Clip shelf base salinity so that it is in the range [4, 40] k/kg. See [@ref HollandJenkins1999].";
    pism_config:ocean.three_equation_model_clip_salinity_option = "clip_shelf_base_salinity";
    pism_config:ocean.three_equation_model_clip_salinity_type = "boolean";

    pism_config:output.backup_interval = 1.0;
    pism_config:output.backup_interval_doc = "wall-clock time between automatic backups";
    pism_config:output.backup_interval_type = "scalar";
    pism_config:output.backup_interval_units = "hours";
    pism_config:output.backup_interval_option = "backup_interval";

    pism_config:output.backup_size = "small";
    pism_config:output.backup_size_choices = "none,small,medium,big_2d,big";
    pism_config:output.backup_size_doc = "The 'size' of a backup file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_config:output.backup_size_option = "backup_size";
    pism_config:output.backup_size_type = "keyword";

    pism_config:output.fill_value = -2e9;
    pism_config:output.fill_value_doc = "_FillValue used when saving diagnostic quantities";
    pism_config:output.fill_value_type = "scalar";
    pism_config:output.fill_value_units = "none";

    pism_config:output.format = "netcdf3";
    pism_config:output.format_choices = "netcdf3,quilt,netcdf4_parallel,pnetcdf";
    pism_config:output.format_doc = "The I/O format used for spatial fields; 'netcdf3' is the default, 'netcd4_parallel' is available if PISM was built with parallel NetCDF-4, and 'pnetcdf' is available if PISM was built with PnetCDF.";
    pism_config:output.format_option = "o_format";
    pism_config:output.format_type = "keyword";

    pism_config:output.ice_free_thickness_standard = 10.0;
    pism_config:output.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a grid cell is considered ice-free for purposes of reporting glacierized area, volume, etc.";
    pism_config:output.ice_free_thickness_standard_type = "scalar";
    pism_config:output.ice_free_thickness_standard_units = "meters";

    pism_config:output.runtime.area_scale_factor_log10 = 6;
    pism_config:output.runtime.area_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for area (in km^2) in summary line to stdout";
    pism_config:output.runtime.area_scale_factor_log10_option = "summary_area_scale_factor_log10";
    pism_config:output.runtime.area_scale_factor_log10_type = "integer";
    pism_config:output.runtime.area_scale_factor_log10_units = "pure number";

    pism_config:output.file_name = "unnamed.nc";
    pism_config:output.file_name_doc = "The file to save final model results to.";
    pism_config:output.file_name_type = "string";
    pism_config:output.file_name_option = "o";

    pism_config:output.runtime.time_unit_name = "year";
    pism_config:output.runtime.time_unit_name_doc = "Time units used when printing model time, time step, and maximum horizontal velocity at summary to stdout.  Must be valid udunits for time.  (E.g. choose from year,month,day,hour,minute,second.)";
    pism_config:output.runtime.time_unit_name_type = "string";

    pism_config:output.runtime.time_use_calendar = "yes";
    pism_config:output.runtime.time_use_calendar_doc = "Whether to use the current calendar when printing model time in summary to stdout.";
    pism_config:output.runtime.time_use_calendar_type = "boolean";

    pism_config:output.runtime.viewer.size = 320;
    pism_config:output.runtime.viewer.size_doc = "default diagnostic viewer size (number of pixels of the longer side)";
    pism_config:output.runtime.viewer.size_option = "view_size";
    pism_config:output.runtime.viewer.size_type = "integer";
    pism_config:output.runtime.viewer.size_units = "count";

    pism_config:output.runtime.viewer.variables = "";
    pism_config:output.runtime.viewer.variables_doc = "comma-separated list of map-plane diagnostic quantities to view at runtime";
    pism_config:output.runtime.viewer.variables_option = "view";
    pism_config:output.runtime.viewer.variables_type = "string";

    pism_config:output.runtime.volume_scale_factor_log10 = 6;
    pism_config:output.runtime.volume_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for volume (in km^3) in summary line to stdout";
    pism_config:output.runtime.volume_scale_factor_log10_option = "summary_vol_scale_factor_log10";
    pism_config:output.runtime.volume_scale_factor_log10_type = "integer";
    pism_config:output.runtime.volume_scale_factor_log10_units = "pure number";

    pism_config:output.save_size = "small";
    pism_config:output.save_size_choices = "none,small,medium,big_2d,big";
    pism_config:output.save_size_doc = "The 'size' of a snapshot file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_config:output.save_size_option = "save_size";
    pism_config:output.save_size_type = "keyword";

    pism_config:output.size = "medium";
    pism_config:output.size_choices = "none,small,medium,big_2d,big";
    pism_config:output.size_doc = "The 'size' of an output file. See configuration parameters output.sizes.medium, output.sizes.big_2d, output.sizes.big";
    pism_config:output.size_option = "o_size";
    pism_config:output.size_type = "keyword";

    pism_config:output.sizes.big = "cts,liqfrac,temp,temp_pa,uvel,vvel,wvel,wvel_rel";
    pism_config:output.sizes.big_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables and variables listed in output.sizes.medium and output.sizes.big_2d) if 'big' output size is selected. Does not include fields written by sub-models.";
    pism_config:output.sizes.big_type = "string";

    pism_config:output.sizes.big_2d = "age,bfrict,bheatflx,bmelt,bwp,bwprel,cell_area,dbdt,effbwp,enthalpybase,enthalpysurf,flux_divergence,hardav,hydroinput,lat,litho_temp,lon,nuH,ocean_kill_mask,rank,tempbase,tempicethk,tempicethk_basal,temppabase,tempsurf,thk,thksmooth,tillphi,topg,velbar,velbase,wallmelt,wvelbase";
    pism_config:output.sizes.big_2d_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables and variables listed in output.sizes.medium) if 'big_2d' output size is selected. Does not include fields written by boundary models.";
    pism_config:output.sizes.big_2d_type = "string";

    pism_config:output.sizes.medium = "bwat,bwatvel,climatic_mass_balance,diffusivity,enthalpy,flux,flux_mag,ice_surface_temp,liqfrac,mask,schoofs_theta,strain_rates,taub_mag,tauc,taud_mag,temp_pa,tillwat,topgsmooth,usurf,velbar_mag,velbase_mag,velsurf,velsurf_mag,wvelsurf";
    pism_config:output.sizes.medium_doc = "Comma-separated list of variables to write to the output (in addition to model_state variables) if 'medium' output size (the default) is selected. Does not include fields written by sub-models.";
    pism_config:output.sizes.medium_type = "string";

    pism_config:output.timeseries.buffer_size = 10000;
    pism_config:output.timeseries.buffer_size_doc = "Number of scalar diagnostic time-series records to hold in memory before writing to disk. (PISM writes this many time-series records to reduce I/O costs.) Send the USR2 signal to flush time-series.";
    pism_config:output.timeseries.buffer_size_type = "integer";
    pism_config:output.timeseries.buffer_size_units = "count";

    pism_config:output.timeseries.variables = "";
    pism_config:output.timeseries.variables_doc = "Requested scalar (time-series) diagnostics. Leave empty to save all available diagnostics.";
    pism_config:output.timeseries.variables_option = "ts_vars";
    pism_config:output.timeseries.variables_type = "string";

    pism_config:output.timeseries.append = "false";
    pism_config:output.timeseries.append_type = "boolean";
    pism_config:output.timeseries.append_option = "ts_append";
    pism_config:output.timeseries.append_doc = "If true, append to the scalar time series output file.";

    pism_config:output.timeseries.filename = "";
    pism_config:output.timeseries.filename_type = "string";
    pism_config:output.timeseries.filename_option = "ts_file";
    pism_config:output.timeseries.filename_doc = "Name of the file to save scalar time series to. Leave empty to disable reporting scalar time-series.";

    pism_config:output.variable_order = "yxz";
    pism_config:output.variable_order_choices = "xyz,yxz,zyx";
    pism_config:output.variable_order_doc = "Variable order to use in output files.";
    pism_config:output.variable_order_option = "o_order";
    pism_config:output.variable_order_type = "keyword";

    pism_config:regional.no_model_strip = 5.0;
    pism_config:regional.no_model_strip_doc = "Default width of the 'no model strip' in regional setups.";
    pism_config:regional.no_model_strip_option = "no_model_strip";
    pism_config:regional.no_model_strip_type = "scalar";
    pism_config:regional.no_model_strip_units = "km";

    pism_config:regional.zero_gradient = "false";
    pism_config:regional.zero_gradient_type = "boolean";
    pism_config:regional.zero_gradient_option = "zero_grad_where_no_model";
    pism_config:regional.zero_gradient_doc = "Use zero ice thickness and ice surface gradient in the no_model_mask area.";

    pism_config:run_info.institution = "";
    pism_config:run_info.institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";
    pism_config:run_info.institution_option = "institution";
    pism_config:run_info.institution_type = "string";

    pism_config:run_info.title = "";
    pism_config:run_info.title_doc = "Free-form string containing a concise description of the current run. This string is written to output files as the 'title' global attribute.";
    pism_config:run_info.title_option = "title";
    pism_config:run_info.title_type = "string";

    pism_config:stress_balance.calving_front_stress_bc = "no";
    pism_config:stress_balance.calving_front_stress_bc_doc = "Apply CFBC condition as in [@ref Albrechtetal2011, @ref Winkelmannetal2011].  May only apply to some stress balances; e.g. SSAFD as of May 2011.  If not set then a strength-extension is used, as in [@ref BBssasliding].";
    pism_config:stress_balance.calving_front_stress_bc_option = "cfbc";
    pism_config:stress_balance.calving_front_stress_bc_type = "boolean";

    pism_config:stress_balance.ice_free_thickness_standard = 10.0;
    pism_config:stress_balance.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a cell is considered ice-free for purposes of computing ice velocity distribution.";
    pism_config:stress_balance.ice_free_thickness_standard_type = "scalar";
    pism_config:stress_balance.ice_free_thickness_standard_units = "meters";

    pism_config:stress_balance.model = "sia";
    pism_config:stress_balance.model_choices = "none,prescribed_sliding,sia,ssa,prescribed_sliding+sia,ssa+sia";
    pism_config:stress_balance.model_doc = "Stress balance model";
    pism_config:stress_balance.model_option = "stress_balance";
    pism_config:stress_balance.model_type = "keyword";

    pism_config:stress_balance.sia.Glen_exponent = 3.0;
    pism_config:stress_balance.sia.Glen_exponent_doc = "Glen exponent in ice flow law for SIA";
    pism_config:stress_balance.sia.Glen_exponent_option = "sia_n";
    pism_config:stress_balance.sia.Glen_exponent_type = "scalar";
    pism_config:stress_balance.sia.Glen_exponent_units = "pure number";

    pism_config:stress_balance.sia.bed_smoother_range = 5.0e3;
    pism_config:stress_balance.sia.bed_smoother_range_doc = "half-width of smoothing domain for stressbalance::BedSmoother, in implementing [@ref Schoofbasaltopg2003] bed roughness parameterization for SIA; set value to zero to turn off mechanism";
    pism_config:stress_balance.sia.bed_smoother_range_option = "bed_smoother_range";
    pism_config:stress_balance.sia.bed_smoother_range_type = "scalar";
    pism_config:stress_balance.sia.bed_smoother_range_units = "meters";

    pism_config:stress_balance.sia.e_age_coupling = "no";
    pism_config:stress_balance.sia.e_age_coupling_doc = "Couple the SIA enhancement factor to age as in [@ref Greve].";
    pism_config:stress_balance.sia.e_age_coupling_option = "e_age_coupling";
    pism_config:stress_balance.sia.e_age_coupling_type = "boolean";

    pism_config:stress_balance.sia.enhancement_factor = 1.0;
    pism_config:stress_balance.sia.enhancement_factor_doc = "Flow enhancement factor for SIA";
    pism_config:stress_balance.sia.enhancement_factor_option = "sia_e";
    pism_config:stress_balance.sia.enhancement_factor_type = "scalar";
    pism_config:stress_balance.sia.enhancement_factor_units = "1";

    pism_config:stress_balance.sia.enhancement_factor_interglacial = 1.0;
    pism_config:stress_balance.sia.enhancement_factor_interglacial_doc = "Flow enhancement factor for SIA; used for ice accumulated during interglacial periods.";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_option = "sia_e_interglacial";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_type = "scalar";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_units = "1";

    pism_config:stress_balance.sia.flow_law = "gpbld";
    pism_config:stress_balance.sia.flow_law_choices = "arr,arrwarm,gk,gpbld,hooke,isothermal_glen,pb,gpbld3";
    pism_config:stress_balance.sia.flow_law_doc = "The SIA flow law.";
    pism_config:stress_balance.sia.flow_law_option = "sia_flow_law";
    pism_config:stress_balance.sia.flow_law_type = "keyword";

    pism_config:stress_balance.sia.grain_size_age_coupling = "no";
    pism_config:stress_balance.sia.grain_size_age_coupling_doc = "Use age of the ice to compute grain size to use with the Goldsby-Kohlstedt [@ref GoldsbyKohlstedt] flow law";
    pism_config:stress_balance.sia.grain_size_age_coupling_option = "grain_size_age_coupling";
    pism_config:stress_balance.sia.grain_size_age_coupling_type = "boolean";

    pism_config:stress_balance.sia.surface_gradient_method = "haseloff";
    pism_config:stress_balance.sia.surface_gradient_method_choices = "eta,haseloff,mahaffy";
    pism_config:stress_balance.sia.surface_gradient_method_doc = "method used for surface gradient calculation at staggered grid points";
    pism_config:stress_balance.sia.surface_gradient_method_option = "gradient";
    pism_config:stress_balance.sia.surface_gradient_method_type = "keyword";

    pism_config:stress_balance.ssa.Glen_exponent = 3.0;
    pism_config:stress_balance.ssa.Glen_exponent_doc = "Glen exponent in ice flow law for SSA";
    pism_config:stress_balance.ssa.Glen_exponent_option = "ssa_n";
    pism_config:stress_balance.ssa.Glen_exponent_type = "scalar";
    pism_config:stress_balance.ssa.Glen_exponent_units = "pure number";

    pism_config:stress_balance.ssa.compute_surface_gradient_inward = "no";
    pism_config:stress_balance.ssa.compute_surface_gradient_inward_doc = "If yes then use inward first-order differencing in computing surface gradient in the SSA objects.";
    pism_config:stress_balance.ssa.compute_surface_gradient_inward_type = "boolean";

    pism_config:stress_balance.ssa.dirichlet_bc = "no";
    pism_config:stress_balance.ssa.dirichlet_bc_doc = "apply SSA velocity Dirichlet boundary condition";
    pism_config:stress_balance.ssa.dirichlet_bc_option = "ssa_dirichlet_bc";
    pism_config:stress_balance.ssa.dirichlet_bc_type = "boolean";

    pism_config:stress_balance.ssa.enhancement_factor = 1.0;
    pism_config:stress_balance.ssa.enhancement_factor_doc = "Flow enhancement factor for SSA";
    pism_config:stress_balance.ssa.enhancement_factor_option = "ssa_e";
    pism_config:stress_balance.ssa.enhancement_factor_type = "scalar";
    pism_config:stress_balance.ssa.enhancement_factor_units = "1";

    pism_config:stress_balance.ssa.enhancement_factor_interglacial = 1.0;
    pism_config:stress_balance.ssa.enhancement_factor_interglacial_doc = "Flow enhancement factor for SSA; used for ice accumulated during interglacial periods.";
    pism_config:stress_balance.ssa.enhancement_factor_interglacial_option = "ssa_e_interglacial";
    pism_config:stress_balance.ssa.enhancement_factor_interglacial_type = "scalar";
    pism_config:stress_balance.ssa.enhancement_factor_interglacial_units = "1";

    pism_config:stress_balance.ssa.epsilon = 1.0e13;
    pism_config:stress_balance.ssa.epsilon_doc = "Initial amount of regularization in computation of product of effective viscosity and thickness (nu * H).  This default value for nu * H comes e.g. from a hardness for the Ross ice shelf (bar B) = 1.9e8 Pa s^(1/3) [@ref MacAyealetal] and a typical strain rate of 0.001 year-1 for the Ross ice shelf, giving nu = (bar B) / (2 * 0.001^(2/3)) = 9.49e+14 Pa s ~~ 30 MPa year, the value in [@ref Ritzetal2001], but with a tiny thickness H of about 1 cm.";
    pism_config:stress_balance.ssa.epsilon_option = "ssa_eps";
    pism_config:stress_balance.ssa.epsilon_type = "scalar";
    pism_config:stress_balance.ssa.epsilon_units = "Pascal second meter";

    pism_config:stress_balance.ssa.fd.brutal_sliding = "false";
    pism_config:stress_balance.ssa.fd.brutal_sliding_doc = "Enhance sliding speed brutally.";
    pism_config:stress_balance.ssa.fd.brutal_sliding_option = "brutal_sliding";
    pism_config:stress_balance.ssa.fd.brutal_sliding_type = "boolean";

    pism_config:stress_balance.ssa.fd.brutal_sliding_scale = 1.0;
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_doc = "Brutal SSA Sliding Scale";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_option = "brutal_sliding_scale";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_type = "scalar";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_units = "1";

    pism_config:stress_balance.ssa.fd.lateral_drag.enabled = "false";
    pism_config:stress_balance.ssa.fd.lateral_drag.enabled_doc = "set viscosity at ice shelf margin next to ice free bedrock as friction parameterization";
    pism_config:stress_balance.ssa.fd.lateral_drag.enabled_type = "boolean";

    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity = 5.0e15;
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_doc = "Staggered Viscosity used as side friction parameterization.";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_option = "nu_bedrock";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_type = "scalar";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_units = "Pascal second";

    pism_config:stress_balance.ssa.fd.max_iterations = 300;
    pism_config:stress_balance.ssa.fd.max_iterations_doc = "Maximum number of iterations for the ice viscosity computation, in the SSAFD object";
    pism_config:stress_balance.ssa.fd.max_iterations_option = "ssa_maxi";
    pism_config:stress_balance.ssa.fd.max_iterations_type = "integer";
    pism_config:stress_balance.ssa.fd.max_iterations_units = "count";

    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation = 0.8;
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_doc = "In event of 'Effective viscosity not converged' failure, use outer iteration rule nuH <- nuH + f (nuH - nuH_old), where f is this parameter.";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_option = "ssafd_nuH_iter_failure_underrelaxation";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_type = "scalar";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_units = "pure number";

    pism_config:stress_balance.ssa.fd.relative_convergence = 1.0e-4;
    pism_config:stress_balance.ssa.fd.relative_convergence_doc = "Relative change tolerance for the effective viscosity in the SSAFD object";
    pism_config:stress_balance.ssa.fd.relative_convergence_option = "ssa_rtol";
    pism_config:stress_balance.ssa.fd.relative_convergence_type = "scalar";
    pism_config:stress_balance.ssa.fd.relative_convergence_units = "1";

    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries = "yes";
    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries_doc = "Replace zero diagonal entries in the SSAFD matrix with basal_resistance.beta_ice_free_bedrock to avoid solver failures.";
    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries_type = "boolean";

    pism_config:stress_balance.ssa.flow_law = "gpbld";
    pism_config:stress_balance.ssa.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb,gpbld3";
    pism_config:stress_balance.ssa.flow_law_doc = "The SSA flow law.";
    pism_config:stress_balance.ssa.flow_law_option = "ssa_flow_law";
    pism_config:stress_balance.ssa.flow_law_type = "keyword";

    pism_config:stress_balance.ssa.method = "fd";
    pism_config:stress_balance.ssa.method_choices = "fd,fem";
    pism_config:stress_balance.ssa.method_doc = "Algorithm for computing the SSA solution.";
    pism_config:stress_balance.ssa.method_option = "ssa_method";
    pism_config:stress_balance.ssa.method_type = "keyword";

    pism_config:stress_balance.ssa.strength_extension.constant_nu = 9.48680701906572e+14;
    pism_config:stress_balance.ssa.strength_extension.constant_nu_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  This value for nu comes from hardness (bar B)=1.9e8 Pa s^(1/3) [@ref MacAyealetal] and a typical strain rate of 0.001 year-1:  nu = (bar B) / (2 * 0.001^(2/3)).  Compare the value of 9.45e14 Pa s = 30 MPa year in [@ref Ritzetal2001].";
    pism_config:stress_balance.ssa.strength_extension.constant_nu_type = "scalar";
    pism_config:stress_balance.ssa.strength_extension.constant_nu_units = "Pascal second";

    pism_config:stress_balance.ssa.strength_extension.min_thickness = 50.0;
    pism_config:stress_balance.ssa.strength_extension.min_thickness_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  At ice thicknesses below this value the product nu*H switches from the normal vertical integral to a constant value.  The geometry itself is not affected by this value.";
    pism_config:stress_balance.ssa.strength_extension.min_thickness_type = "scalar";
    pism_config:stress_balance.ssa.strength_extension.min_thickness_units = "meters";

    pism_config:stress_balance.vertical_velocity_approximation = "centered";
    pism_config:stress_balance.vertical_velocity_approximation_choices = "centered,upstream";
    pism_config:stress_balance.vertical_velocity_approximation_doc = "Vertical velocity FD approximation. \"Upstream\" uses first-order finite difference to compute u_x and v_y. Uses basal velocity to make decisions.";
    pism_config:stress_balance.vertical_velocity_approximation_option = "vertical_velocity_approximation";
    pism_config:stress_balance.vertical_velocity_approximation_type = "keyword";

    pism_config:surface.force_to_thickness.alpha = 0.01;
    pism_config:surface.force_to_thickness.alpha_doc = "exponential coefficient in force-to-thickness mechanism";
    pism_config:surface.force_to_thickness.alpha_type = "scalar";
    pism_config:surface.force_to_thickness.alpha_units = "year-1";

    pism_config:surface.force_to_thickness.ice_free_alpha_factor = 1.0;
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_doc = "surface.force_to_thickness.alpha is multiplied by this factor in areas that are ice-free according to the target ice thickness and surface.force_to_thickness.ice_free_thickness_threshold";
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_type = "scalar";
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_units = "1";

    pism_config:surface.force_to_thickness.ice_free_thickness_threshold = 1.0;
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_doc = "threshold of ice thickness in the force-to-thickness target field. Used to determine whether to use surface.force_to_thickness.ice_free_alpha_factor.";
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_type = "scalar";
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_units = "meters";

    pism_config:surface.force_to_thickness.start_time = -4.54e9;
    pism_config:surface.force_to_thickness.start_time_doc = "Starting time for the \"force to thickness\" modifier; the default is \"start from the creation of the Earth.\"";
    pism_config:surface.force_to_thickness.start_time_type = "scalar";
    pism_config:surface.force_to_thickness.start_time_units = "years";

    pism_config:surface.pdd.air_temp_all_precip_as_rain = 275.15;
    pism_config:surface.pdd.air_temp_all_precip_as_rain_doc = "threshold temperature above which all precipitation is rain; must exceed surface.pdd.air_temp_all_precip_as_snow to avoid division by zero, because difference is in a denominator";
    pism_config:surface.pdd.air_temp_all_precip_as_rain_type = "scalar";
    pism_config:surface.pdd.air_temp_all_precip_as_rain_units = "Kelvin";

    pism_config:surface.pdd.air_temp_all_precip_as_snow = 273.15;
    pism_config:surface.pdd.air_temp_all_precip_as_snow_doc = "threshold temperature below which all precipitation is snow";
    pism_config:surface.pdd.air_temp_all_precip_as_snow_type = "scalar";
    pism_config:surface.pdd.air_temp_all_precip_as_snow_units = "Kelvin";

    pism_config:surface.pdd.balance_year_start_day = 274;
    pism_config:surface.pdd.balance_year_start_day_doc = "day of year for October 1st, beginning of the balance year in northern latitudes.";
    pism_config:surface.pdd.balance_year_start_day_type = "integer";
    pism_config:surface.pdd.balance_year_start_day_units = "ordinal day number";

    pism_config:surface.pdd.aschwanden.beta_ice_c = 0.006;
    pism_config:surface.pdd.aschwanden.beta_ice_c_doc = "water-equivalent thickness; for formula (6) in [@ref Aschwandenetal2009] ";
    pism_config:surface.pdd.aschwanden.beta_ice_c_type = "scalar";
    pism_config:surface.pdd.aschwanden.beta_ice_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.aschwanden.beta_ice_w = 0.008;
    pism_config:surface.pdd.aschwanden.beta_ice_w_doc = "water-equivalent thickness; for formula (6) in [@ref Aschwandenetal2009] ";
    pism_config:surface.pdd.aschwanden.beta_ice_w_type = "scalar";
    pism_config:surface.pdd.aschwanden.beta_ice_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.aschwanden.beta_snow_c = 0.0015;
    pism_config:surface.pdd.aschwanden.beta_snow_c_doc = "water-equivalent thickness; for formula (6) in [@ref Aschwandenetal2009] ";
    pism_config:surface.pdd.aschwanden.beta_snow_c_type = "scalar";
    pism_config:surface.pdd.aschwanden.beta_snow_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.aschwanden.beta_snow_w = 0.003;
    pism_config:surface.pdd.aschwanden.beta_snow_w_doc = "water-equivalent thickness; for formula (6) in [@ref Aschwandenetal2009] ";
    pism_config:surface.pdd.aschwanden.beta_snow_w_type = "scalar";
    pism_config:surface.pdd.aschwanden.beta_snow_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.aschwanden.latitude_beta_w = 77.0;
    pism_config:surface.pdd.aschwanden.latitude_beta_w_doc = "latitude below which to use warm case, in formula (6) in [@ref Aschwandenetal2009] ";
    pism_config:surface.pdd.aschwanden.latitude_beta_w_type = "scalar";
    pism_config:surface.pdd.aschwanden.latitude_beta_w_units = "degree_north";

    pism_config:surface.pdd.aschwanden.warm_cold_transition_width = 1.0;
    pism_config:surface.pdd.aschwanden.warm_cold_transition_width_doc = "smoothing width in degrees for linear transition between warm and cold values";
    pism_config:surface.pdd.aschwanden.warm_cold_transition_width_type = "scalar";
    pism_config:surface.pdd.aschwanden.warm_cold_transition_width_units = "degree_north";

    pism_config:surface.pdd.factor_ice = 0.00879120879120879;
    pism_config:surface.pdd.factor_ice_doc = "EISMINT-Greenland value [@ref RitzEISMINT]; = (8 mm liquid-water-equivalent) / (pos degree day)";
    pism_config:surface.pdd.factor_ice_type = "scalar";
    pism_config:surface.pdd.factor_ice_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.factor_snow = 0.0032967032967033;
    pism_config:surface.pdd.factor_snow_doc = "EISMINT-Greenland value [@ref RitzEISMINT]; = (3 mm liquid-water-equivalent) / (pos degree day)";
    pism_config:surface.pdd.factor_snow_type = "scalar";
    pism_config:surface.pdd.factor_snow_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.T_c = 272.15;
    pism_config:surface.pdd.fausto.T_c_doc = "= -1 + 273.15; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.T_c_type = "scalar";
    pism_config:surface.pdd.fausto.T_c_units = "Kelvin";

    pism_config:surface.pdd.fausto.T_w = 283.15;
    pism_config:surface.pdd.fausto.T_w_doc = "= 10 + 273.15; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.T_w_type = "scalar";
    pism_config:surface.pdd.fausto.T_w_units = "Kelvin";

    pism_config:surface.pdd.fausto.beta_ice_c = 0.015;
    pism_config:surface.pdd.fausto.beta_ice_c_doc = "water-equivalent thickness; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.beta_ice_c_type = "scalar";
    pism_config:surface.pdd.fausto.beta_ice_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_ice_w = 0.007;
    pism_config:surface.pdd.fausto.beta_ice_w_doc = "water-equivalent thickness; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.beta_ice_w_type = "scalar";
    pism_config:surface.pdd.fausto.beta_ice_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_snow_c = 0.003;
    pism_config:surface.pdd.fausto.beta_snow_c_doc = "water-equivalent thickness; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.beta_snow_c_type = "scalar";
    pism_config:surface.pdd.fausto.beta_snow_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_snow_w = 0.003;
    pism_config:surface.pdd.fausto.beta_snow_w_doc = "water-equivalent thickness; for formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.beta_snow_w_type = "scalar";
    pism_config:surface.pdd.fausto.beta_snow_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.latitude_beta_w = 72.0;
    pism_config:surface.pdd.fausto.latitude_beta_w_doc = "latitude below which to use warm case, in formula (6) in [@ref Faustoetal2009] ";
    pism_config:surface.pdd.fausto.latitude_beta_w_type = "scalar";
    pism_config:surface.pdd.fausto.latitude_beta_w_units = "degree_north";

    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio = 0.75;
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_doc = "How much firn as a fraction of accumulation is turned into ice";
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_type = "scalar";
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_units = "1";

    pism_config:surface.pdd.firn_depth_file = "";
    pism_config:surface.pdd.firn_depth_file_option = "pdd_firn_depth_file";
    pism_config:surface.pdd.firn_depth_file_doc = "The name of the file to read the firn_depth from.";
    pism_config:surface.pdd.firn_depth_file_type = "string";

    pism_config:surface.pdd.temperature_standard_deviation_file = "";
    pism_config:surface.pdd.temperature_standard_deviation_file_option = "pdd_sd_file";
    pism_config:surface.pdd.temperature_standard_deviation_file_doc = "The name of the file to read air_temp_sd from.";
    pism_config:surface.pdd.temperature_standard_deviation_file_type = "string";

    pism_config:surface.pdd.interpret_precip_as_snow = "no";
    pism_config:surface.pdd.interpret_precip_as_snow_doc = "Interpret precipitation as snow fall.";
    pism_config:surface.pdd.interpret_precip_as_snow_type = "boolean";

    pism_config:surface.pdd.max_evals_per_year = 52;
    pism_config:surface.pdd.max_evals_per_year_doc = "maximum number of times the PDD scheme will ask for air temperature and precipitation to build location-dependent time series for computing (expected) number of positive degree days and snow accumulation; the default means the PDD uses weekly samples of the annual cycle; see also surface.pdd.std_dev";
    pism_config:surface.pdd.max_evals_per_year_type = "integer";
    pism_config:surface.pdd.max_evals_per_year_units = "count";

    pism_config:surface.pdd.positive_threshold_temp = 273.15;
    pism_config:surface.pdd.positive_threshold_temp_doc = "temperature used to determine meaning of 'positive' degree day";
    pism_config:surface.pdd.positive_threshold_temp_type = "scalar";
    pism_config:surface.pdd.positive_threshold_temp_units = "Kelvin";

    pism_config:surface.pdd.refreeze = 0.6;
    pism_config:surface.pdd.refreeze_doc = "EISMINT-Greenland value [@ref RitzEISMINT]";
    pism_config:surface.pdd.refreeze_type = "scalar";
    pism_config:surface.pdd.refreeze_units = "1";

    pism_config:surface.pdd.refreeze_ice_melt = "yes";
    pism_config:surface.pdd.refreeze_ice_melt_doc = "If set to 'yes', refreeze surface.pdd.refreeze fraction of melted ice, otherwise all of the melted ice runs off.";
    pism_config:surface.pdd.refreeze_ice_melt_type = "boolean";

    pism_config:surface.pdd.std_dev = 5.0;
    pism_config:surface.pdd.std_dev_doc = "std dev of daily temp variation; = EISMINT-Greenland value [@ref RitzEISMINT] ";
    pism_config:surface.pdd.std_dev_type = "scalar";
    pism_config:surface.pdd.std_dev_units = "Kelvin";

    pism_config:surface.pdd.std_dev_lapse_lat_base = 72.0;
    pism_config:surface.pdd.std_dev_lapse_lat_base_doc = "std_dev is a function of latitude, with value surface.pdd.std_dev at this latitude; this value only active if surface.pdd.std_dev_lapse_lat_rate is nonzero ";
    pism_config:surface.pdd.std_dev_lapse_lat_base_type = "scalar";
    pism_config:surface.pdd.std_dev_lapse_lat_base_units = "degree_north";

    pism_config:surface.pdd.std_dev_lapse_lat_rate = 0.0;
    pism_config:surface.pdd.std_dev_lapse_lat_rate_doc = "std_dev is a function of latitude, with rate of change with respect to latitude given by this constant ";
    pism_config:surface.pdd.std_dev_lapse_lat_rate_type = "scalar";
    pism_config:surface.pdd.std_dev_lapse_lat_rate_units = "Kelvin / degree_north";

    pism_config:surface.pdd.std_dev_param_a = -0.15;
    pism_config:surface.pdd.std_dev_param_a_doc = "Parameter a in Sigma = a*T + b, with T in degrees C. Used only if surface.pdd.std_dev_use_param is set to yes.";
    pism_config:surface.pdd.std_dev_param_a_type = "scalar";
    pism_config:surface.pdd.std_dev_param_a_units = "pure number";

    pism_config:surface.pdd.std_dev_param_b = 0.66;
    pism_config:surface.pdd.std_dev_param_b_doc = "Parameter b in Sigma = a*T + b, with T in degrees C. Used only if surface.pdd.std_dev_use_param is set to yes.";
    pism_config:surface.pdd.std_dev_param_b_type = "scalar";
    pism_config:surface.pdd.std_dev_param_b_units = "Kelvin";

    pism_config:surface.pdd.std_dev_use_param = "no";
    pism_config:surface.pdd.std_dev_use_param_doc = "Parameterize standard deviation as a linear function of air temperature over ice-covered grid cells. The region of application is controlled by geometry.ice_free_thickness_standard.";
    pism_config:surface.pdd.std_dev_use_param_type = "boolean";

    pism_config:surface.pressure = 0.0;
    pism_config:surface.pressure_doc = "atmospheric pressure; = pressure at ice surface";
    pism_config:surface.pressure_type = "scalar";
    pism_config:surface.pressure_units = "Pascal";

    pism_config:surface.temp_to_runoff_a = 0.5;
    pism_config:surface.temp_to_runoff_a_doc = "a in runoff=a * temp + b";
    pism_config:surface.temp_to_runoff_a_type = "scalar";
    pism_config:surface.temp_to_runoff_a_units = "K-1";

    pism_config:time.calendar = "365_day";
    pism_config:time.calendar_choices = "standard,gregorian,proleptic_gregorian,noleap,365_day,360_day,julian,none";
    pism_config:time.calendar_doc = "The calendar to use.";
    pism_config:time.calendar_option = "calendar";
    pism_config:time.calendar_type = "keyword";

    pism_config:time.dimension_name = "time";
    pism_config:time.dimension_name_doc = "The name of the time dimension in PISM output files.";
    pism_config:time.dimension_name_type = "string";

    pism_config:time.eemian_end = -114500.0;
    pism_config:time.eemian_end_doc = "End of the Eemian interglacial period. See [@ref Greve97Greenland].";
    pism_config:time.eemian_end_type = "scalar";
    pism_config:time.eemian_end_units = "years";

    pism_config:time.eemian_start = -132000.0;
    pism_config:time.eemian_start_doc = "Start of the Eemian interglacial period. See [@ref Greve97Greenland].";
    pism_config:time.eemian_start_type = "scalar";
    pism_config:time.eemian_start_units = "years";

    pism_config:time.holocene_start = -11000.0;
    pism_config:time.holocene_start_doc = "Start of the Holocene interglacial period. See [@ref Greve97Greenland].";
    pism_config:time.holocene_start_type = "scalar";
    pism_config:time.holocene_start_units = "years";

    pism_config:time.reference_date = "1-1-1";
    pism_config:time.reference_date_doc = "year-month-day; reference date used for calendar computations and in PISM output files";
    pism_config:time.reference_date_type = "string";

    pism_config:time.run_length = 1000;
    pism_config:time.run_length_doc = "Default run length";
    pism_config:time.run_length_type = "scalar";
    pism_config:time.run_length_units = "years";

    pism_config:time.start_year = 0;
    pism_config:time.start_year_doc = "Start year.";
    pism_config:time.start_year_type = "scalar";
    pism_config:time.start_year_units = "years";

    pism_config:time_stepping.adaptive_ratio = 0.12;
    pism_config:time_stepping.adaptive_ratio_doc = "Adaptive time stepping ratio for the explicit scheme for the mass balance equation; @ref BBL, inequality (25)";
    pism_config:time_stepping.adaptive_ratio_option = "adapt_ratio";
    pism_config:time_stepping.adaptive_ratio_type = "scalar";
    pism_config:time_stepping.adaptive_ratio_units = "1";

    pism_config:time_stepping.count_steps = "no";
    pism_config:time_stepping.count_steps_doc = "If yes, IceModel::run() will count the number of time steps it took.  Sometimes useful for performance evaluation.  Counts all steps, regardless of whether processes (mass continuity, energy, velocity, ...) occurred within the step.";
    pism_config:time_stepping.count_steps_option = "count_steps";
    pism_config:time_stepping.count_steps_type = "boolean";

    pism_config:time_stepping.hit_extra_times = "yes";
    pism_config:time_stepping.hit_extra_times_doc = "Modify the time-stepping mechanism to hit times requested using -extra_times.";
    pism_config:time_stepping.hit_extra_times_option = "extra_force_output_times";
    pism_config:time_stepping.hit_extra_times_type = "boolean";

    pism_config:time_stepping.hit_multiples = 0.0;
    pism_config:time_stepping.hit_multiples_doc = "Hit every X years, where X is specified using this parameter. Use 0 to disable";
    pism_config:time_stepping.hit_multiples_option = "timestep_hit_multiples";
    pism_config:time_stepping.hit_multiples_type = "scalar";
    pism_config:time_stepping.hit_multiples_units = "years";

    pism_config:time_stepping.hit_save_times = "no";
    pism_config:time_stepping.hit_save_times_doc = "Modify the time-stepping mechanism to hit times requested using -save_times.";
    pism_config:time_stepping.hit_save_times_option = "save_force_output_times";
    pism_config:time_stepping.hit_save_times_type = "boolean";

    pism_config:time_stepping.hit_ts_times = "no";
    pism_config:time_stepping.hit_ts_times_doc = "Modify the time-stepping mechanism to hit times requested using -ts_times.";
    pism_config:time_stepping.hit_ts_times_type = "boolean";

    pism_config:time_stepping.maximum_time_step = 60.0;
    pism_config:time_stepping.maximum_time_step_doc = "Maximum allowed time step length";
    pism_config:time_stepping.maximum_time_step_option = "max_dt";
    pism_config:time_stepping.maximum_time_step_type = "scalar";
    pism_config:time_stepping.maximum_time_step_units = "years";

    pism_config:time_stepping.skip.enabled = "no";
    pism_config:time_stepping.skip.enabled_doc = "Use the temperature, age, and SSA stress balance computation skipping mechanism.";
    pism_config:time_stepping.skip.enabled_option = "skip";
    pism_config:time_stepping.skip.enabled_type = "boolean";

    pism_config:time_stepping.skip.max = 10;
    pism_config:time_stepping.skip.max_doc = "Number of mass-balance steps, including SIA diffusivity updates, to perform before a the temperature, age, and SSA stress balance computations are done";
    pism_config:time_stepping.skip.max_option = "skip_max";
    pism_config:time_stepping.skip.max_type = "integer";
    pism_config:time_stepping.skip.max_units = "count";

    pism_config:long_name = "PISM configuration flags and parameters.";
    pism_config:long_name_doc = "The 'long_name' attribute is required by CF conventions. It is not used by PISM itself.";
}
