netcdf grid {
dimensions:
// length of the x dimension is not important
  x = 1 ;
// length of the y dimension is not important
  y = 1 ;
  nv2 = 2 ;
variables:
  double x(x) ;
    x:units = "m" ;
    x:standard_name = "projection_x_coordinate" ;
    x:bounds = "x_bnds";
  double x_bnds(x, nv2);
  double y(y) ;
    y:units = "m" ;
    y:standard_name = "projection_y_coordinate" ;
    y:bounds = "y_bnds";
  double y_bnds(y, nv2);
  byte domain;
    domain:dimensions = "x y";
    domain:grid_mapping = "mapping";
  byte mapping;
    mapping:proj_params = "EPSG:3413";

// global attributes:
  :Conventions = "CF-1.11";

data:
// x values are not used
   x = 100000.0 ;
   x_bnds = -800000.0, 1000000.0;
// x values are not used
   y = -1997500.0 ;
   y_bnds = -3400000, -595000;
}
