// Copyright (C) 2007--2008 Jed Brown and Ed Bueler
//
// This file is part of PISM.
//
// PISM is free software; you can redistribute it and/or modify it under the
// terms of the GNU General Public License as published by the Free Software
// Foundation; either version 2 of the License, or (at your option) any later
// version.
//
// PISM is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS
// FOR A PARTICULAR PURPOSE.  See the GNU General Public License for more
// details.
//
// You should have received a copy of the GNU General Public License
// along with PISM; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA  02110-1301  USA


// regarding attribute "pism_intent": pism_intent can have one of five values:
//           model_state, mapping, climate_steady, climate_snapshot, diagnostic
//
// 1.  those variables with pism_intent attribute "model_state" are *required* if the .nc file is
//     to be used to initialize PISM (by "-if", i.e. without bootstrapping)
// 2.  those variables with "mapping" are not model state but are generally required by PISM and generally
//     will affect programs which display or process nc files
// 3.  those variables with "climate_steady" or "climate_snapshot" are boundary
//     conditions stored from an earlier bootstrap, or are initialized to constants, but these could be 
//     variables modified by external models (e.g. of ocean or atmosphere ...); modifying these variables 
//     will usually effect the behavior of the PISM run from "-if"
// 4.  "climate_steady" means that the run occurred from bootstrapping information that had no time dimension
//     or had only one time value, and that this variable did not change during the run; "climate_snapshot"
//     otherwise (i.e. -forcing was used or that there was climate data fed from another model)
// 5.  pism_intent "diagnostic" means just that; modifying or removing them will have no effect
//     on the future run

netcdf pism_state { // name is magic in ncgen.rb

dimensions:
  x = 91; // numbers are magic in ncgen.rb
  y = 92;
  z = 93;
  zb = 94;
  t = UNLIMITED;

variables: // The names of variables are magic in PISM source.
  int polar_stereographic;  
    // the following choices are clearly tied to Antarctic but they are only defaults because
    // if the input or bootstrap file has this var then it is written into the pism state file
    polar_stereographic:grid_mapping_name = "polar_stereographic";
    polar_stereographic:straight_vertical_longitude_from_pole = 0.0;
    polar_stereographic:latitude_of_projection_origin = -90.0;
    polar_stereographic:standard_parallel = -71.0;
    polar_stereographic:pism_intent = "mapping";
  // note accuracy desirable for the locations of the points of the grid
  // accuracy is desirable for t(t) even for long runs (e.g. day accuracy for 1e6 year runs
  // so that PDD method works; also note appearance of year at each restart)
  double x(x);
    x:axis = "X";
    x:long_name = "x-coordinate in Cartesian system";
    x:standard_name = "projection_x_coordinate";
    x:units = "m";
    x:pism_intent = "mapping";
  double y(y);
    y:axis = "Y";
    y:long_name = "y-coordinate in Cartesian system";
    y:standard_name = "projection_y_coordinate";
    y:units = "m";
    y:pism_intent = "mapping";
  double z(z);
    z:axis = "Z";
    z:long_name = "z-coordinate in Cartesian system";
    z:standard_name = "projection_z_coordinate";
    z:units = "m";
    z:positive = "up";
    z:pism_intent = "mapping";
  double zb(zb);
    zb:long_name = "z-coordinate in bedrock";
    zb:standard_name = "projection_z_coordinate_in_bedrock";
    zb:units = "m";
    zb:positive = "up";
    zb:pism_intent = "mapping";
  double t(t);
    t:long_name = "time";
    t:units = "seconds since 2007-01-01 00:00:00";
    t:calendar = "none";
    t:axis = "T";
  float lon(t,x,y);
    lon:long_name = "longitude";
    lon:standard_name = "longitude";
    lon:units = "degrees_east";
    lon:pism_intent = "mapping";
  float lat(t,x,y);
    lat:long_name = "latitude";
    lat:standard_name = "latitude";
    lat:units = "degrees_north";
    lat:pism_intent = "mapping";

// 2-dimensional integer mask
  byte mask(t,x,y);
    mask:long_name = "grounded_dragging_floating integer mask";
    mask:pism_intent = "model_state";

// 2-dimensional model quantities
  float thk(t,x,y);
    thk:long_name = "land ice thickness";
    thk:standard_name = "land_ice_thickness";
    thk:units = "m";
    thk:pism_intent = "model_state";
  float bwat(t,x,y);
    bwat:long_name = "effective thickness of subglacial melt water";
    bwat:units = "m";
    bwat:pism_intent = "model_state";
  float topg(t,x,y);
    topg:long_name = "bedrock surface elevation";
    topg:standard_name = "bedrock_altitude";
    topg:units = "m";
    topg:pism_intent = "model_state";
  float dbdt(t,x,y);
    dbdt:long_name = "bedrock uplift rate";
    dbdt:standard_name = "tendency_of_bedrock_altitude";
    dbdt:units = "m s-1";
    dbdt:pism_intent = "model_state";  // note LC bed model treats as model state

// 3-dimensional model quantities
  float temp(t,x,y,z);
    temp:long_name = "ice temperature";
    temp:standard_name = "land_ice_temperature";
    temp:units = "K";
    temp:pism_intent = "model_state";
  float litho_temp(t,x,y,zb);
    litho_temp:long_name = "bedrock temperature";
    litho_temp:standard_name = "bedrock_temperature";
    litho_temp:units = "K";
    litho_temp:pism_intent = "model_state";
  float age(t,x,y,z);
    age:long_name = "age of ice";
    age:standard_name = "land_ice_age";
    age:units = "s";
    age:pism_intent = "model_state";

// 2-dimensional climate or boundary quantities
  float artm(t,x,y);
    artm:long_name = "annual mean air temperature at ice surface";
    artm:standard_name = "surface_temperature";
    artm:units = "K";
    artm:pism_intent = "climate_steady";  // at this point; change to default "climate_snapshot" according
                                        // to -forcing?
  float bheatflx(t,x,y);
    bheatflx:long_name = "upward geothermal flux at bedrock surface";
    bheatflx:units = "W m-2";
    bheatflx:pism_intent = "climate_steady";  // at this point; ditto
  float acab(t,x,y);
    acab:long_name = "mean annual net ice equivalent accumulation (ablation) rate";
    acab:standard_name = "land_ice_surface_specific_mass_balance";
    acab:units = "m s-1";
    acab:pism_intent = "climate_steady";  // at this point; ditto
  float tillphi(t,x,y);
    tillphi:long_name = "friction angle for till under grounded ice sheet";
    tillphi:units = "degrees";
    tillphi:pism_intent = "climate_steady";

// 2-dimensional diagnostic quantities
  float usurf(t,x,y);
    usurf:long_name = "ice upper surface elevation";
    usurf:standard_name = "surface_altitude";
    usurf:units = "m";
    usurf:pism_intent = "diagnostic";  // because h = H + b; H and b are model_state
  float dHdt(t,x,y);
    dHdt:long_name = "rate of change of ice thickness";
    dHdt:units = "m year-1";
    dHdt:pism_intent = "diagnostic";
  float cbar(t,x,y);
    cbar:long_name = "magnitude of vertically-integrated horizontal velocity of ice";
    cbar:units = "m year-1";
    cbar:pism_intent = "diagnostic";
  float cbase(t,x,y);
    cbase:long_name = "magnitude of horizontal velocity of ice at base of ice";
    cbase:units = "m year-1";
    cbase:pism_intent = "diagnostic";
  float csurf(t,x,y);
    csurf:long_name = "magnitude of horizontal velocity of ice at ice surface";
    csurf:units = "m year-1";
    csurf:pism_intent = "diagnostic";
  float wsurf(t,x,y);
    wsurf:long_name = "vertical velocity of ice at ice surface";
    wsurf:units = "m year-1";
    wsurf:pism_intent = "diagnostic";
  float cflx(t,x,y);
    cflx:long_name = "magnitude of vertically-integrated horizontal flux of ice";
    cflx:units = "m2 year-1";
    cflx:pism_intent = "diagnostic";
  float taub(t,x,y);
    taub:long_name = "magnitude of driving shear stress at base of ice";
    taub:units = "Pa";  // Pascals; 100 kPa = 1e5 Pa = 1 bar
    taub:pism_intent = "diagnostic";
  float tauc(t,x,y);
    tauc:long_name = "yield stress for basal till (plastic or pseudo-plastic model)";
    tauc:units = "Pa";  // Pascals; 100 kPa = 1e5 Pa = 1 bar
    tauc:pism_intent = "diagnostic";

// global attributes
    :Conventions = "CF-1.0";

}
