netcdf pism_config {
    variables:
    byte pism_config;

    pism_config:age.enabled = "no";
    pism_config:age.enabled_doc = "Solve age equation (advection equation for ice age).";
    pism_config:age.enabled_option = "age";
    pism_config:age.enabled_type = "flag";

    pism_config:age.initial_value = 0.0;
    pism_config:age.initial_value_doc = "Initial age of ice";
    pism_config:age.initial_value_type = "number";
    pism_config:age.initial_value_units = "years";

    pism_config:atmosphere.anomaly.file = "";
    pism_config:atmosphere.anomaly.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:atmosphere.anomaly.file_option = "atmosphere_anomaly_file";
    pism_config:atmosphere.anomaly.file_type = "string";

    pism_config:atmosphere.anomaly.periodic = "no";
    pism_config:atmosphere.anomaly.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.anomaly.periodic_type = "flag";

    pism_config:atmosphere.delta_P.file = "";
    pism_config:atmosphere.delta_P.file_doc = "Name of the file containing scalar precipitation offsets.";
    pism_config:atmosphere.delta_P.file_option = "atmosphere_delta_P_file";
    pism_config:atmosphere.delta_P.file_type = "string";

    pism_config:atmosphere.delta_P.periodic = "no";
    pism_config:atmosphere.delta_P.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.delta_P.periodic_type = "flag";

    pism_config:atmosphere.delta_T.file = "";
    pism_config:atmosphere.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_config:atmosphere.delta_T.file_option = "atmosphere_delta_T_file";
    pism_config:atmosphere.delta_T.file_type = "string";

    pism_config:atmosphere.delta_T.periodic = "no";
    pism_config:atmosphere.delta_T.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.delta_T.periodic_type = "flag";

    pism_config:atmosphere.elevation_change.file = "";
    pism_config:atmosphere.elevation_change.file_doc = "Name of the file containing the reference surface elevation field (variable :var:`usurf`).";
    pism_config:atmosphere.elevation_change.file_option = "atmosphere_lapse_rate_file";
    pism_config:atmosphere.elevation_change.file_type = "string";

    pism_config:atmosphere.elevation_change.periodic = "no";
    pism_config:atmosphere.elevation_change.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.elevation_change.periodic_type = "flag";

    pism_config:atmosphere.elevation_change.precipitation.lapse_rate = 0.0;
    pism_config:atmosphere.elevation_change.precipitation.lapse_rate_doc = "Elevation lapse rate for the precipitation";
    pism_config:atmosphere.elevation_change.precipitation.lapse_rate_option = "precip_lapse_rate";
    pism_config:atmosphere.elevation_change.precipitation.lapse_rate_type = "number";
    pism_config:atmosphere.elevation_change.precipitation.lapse_rate_units = "(kg m-2 / year) / km";

    pism_config:atmosphere.elevation_change.precipitation.method = "shift";
    pism_config:atmosphere.elevation_change.precipitation.method_choices = "scale,shift";
    pism_config:atmosphere.elevation_change.precipitation.method_doc = "Choose the precipitation adjustment method. ``scale``: use temperature-change-dependent scaling factor. ``shift``: use the precipitation lapse rate.";
    pism_config:atmosphere.elevation_change.precipitation.method_option = "precip_adjustment";
    pism_config:atmosphere.elevation_change.precipitation.method_type = "keyword";

    pism_config:atmosphere.elevation_change.precipitation.temp_lapse_rate = 0.0;
    pism_config:atmosphere.elevation_change.precipitation.temp_lapse_rate_doc = "Elevation lapse rate for the surface temperature used to compute `\\Delta T` in the precipitation scaling factor `\\exp(C \\cdot \\Delta T)`";
    pism_config:atmosphere.elevation_change.precipitation.temp_lapse_rate_option = "precip_temp_lapse_rate";
    pism_config:atmosphere.elevation_change.precipitation.temp_lapse_rate_type = "number";
    pism_config:atmosphere.elevation_change.precipitation.temp_lapse_rate_units = "Kelvin / km";

    pism_config:atmosphere.elevation_change.temperature_lapse_rate = 0.0;
    pism_config:atmosphere.elevation_change.temperature_lapse_rate_doc = "Elevation lapse rate for the surface temperature";
    pism_config:atmosphere.elevation_change.temperature_lapse_rate_option = "temp_lapse_rate";
    pism_config:atmosphere.elevation_change.temperature_lapse_rate_type = "number";
    pism_config:atmosphere.elevation_change.temperature_lapse_rate_units = "Kelvin / km";

    pism_config:atmosphere.fausto_air_temp.c_ma = -0.7189;
    pism_config:atmosphere.fausto_air_temp.c_ma_doc = "latitude-dependence coefficient for formula (1) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.c_ma_type = "number";
    pism_config:atmosphere.fausto_air_temp.c_ma_units = "Kelvin / degree_north";

    pism_config:atmosphere.fausto_air_temp.c_mj = -0.1585;
    pism_config:atmosphere.fausto_air_temp.c_mj_doc = "latitude-dependence coefficient for formula (2) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.c_mj_type = "number";
    pism_config:atmosphere.fausto_air_temp.c_mj_units = "Kelvin / degree_north";

    pism_config:atmosphere.fausto_air_temp.d_ma = 314.98;
    pism_config:atmosphere.fausto_air_temp.d_ma_doc = "41.83+273.15; base temperature for formula (1) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.d_ma_type = "number";
    pism_config:atmosphere.fausto_air_temp.d_ma_units = "Kelvin";

    pism_config:atmosphere.fausto_air_temp.d_mj = 287.85;
    pism_config:atmosphere.fausto_air_temp.d_mj_doc = "= 14.70+273.15; base temperature for formula (2) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.d_mj_type = "number";
    pism_config:atmosphere.fausto_air_temp.d_mj_units = "Kelvin";

    pism_config:atmosphere.fausto_air_temp.gamma_ma = -0.006309;
    pism_config:atmosphere.fausto_air_temp.gamma_ma_doc = "= -6.309 / 1km; mean slope lapse rate for formula (1) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.gamma_ma_type = "number";
    pism_config:atmosphere.fausto_air_temp.gamma_ma_units = "Kelvin / meter";

    pism_config:atmosphere.fausto_air_temp.gamma_mj = -0.005426;
    pism_config:atmosphere.fausto_air_temp.gamma_mj_doc = "= -5.426 / 1km; mean slope lapse rate for formula (2) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.gamma_mj_type = "number";
    pism_config:atmosphere.fausto_air_temp.gamma_mj_units = "Kelvin / meter";

    pism_config:atmosphere.fausto_air_temp.kappa_ma = 0.0672;
    pism_config:atmosphere.fausto_air_temp.kappa_ma_doc = "longitude-dependence coefficient for formula (1) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.kappa_ma_type = "number";
    pism_config:atmosphere.fausto_air_temp.kappa_ma_units = "Kelvin / degree_west";

    pism_config:atmosphere.fausto_air_temp.kappa_mj = 0.0518;
    pism_config:atmosphere.fausto_air_temp.kappa_mj_doc = "longitude-dependence coefficient for formula (2) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.kappa_mj_type = "number";
    pism_config:atmosphere.fausto_air_temp.kappa_mj_units = "Kelvin / degree_west";

    pism_config:atmosphere.fausto_air_temp.summer_peak_day = 196;
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_doc = "day of year for July 15; used in corrected formula (4) in :cite:`Faustoetal2009`";
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_type = "integer";
    pism_config:atmosphere.fausto_air_temp.summer_peak_day_units = "ordinal day number";

    pism_config:atmosphere.frac_P.file = "";
    pism_config:atmosphere.frac_P.file_doc = "Name of the file containing scalar precipitation scaling.";
    pism_config:atmosphere.frac_P.file_option = "atmosphere_frac_P_file";
    pism_config:atmosphere.frac_P.file_type = "string";

    pism_config:atmosphere.frac_P.periodic = "no";
    pism_config:atmosphere.frac_P.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.frac_P.periodic_type = "flag";

    pism_config:atmosphere.given.air_temperature_interpolation = "piecewise_linear";
    pism_config:atmosphere.given.air_temperature_interpolation_choices = "piecewise_linear,piecewise_constant";
    pism_config:atmosphere.given.air_temperature_interpolation_doc = "Temporal interpolation type used for near-surface air temperatures";
    pism_config:atmosphere.given.air_temperature_interpolation_type = "keyword";

    pism_config:atmosphere.given.file = "";
    pism_config:atmosphere.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:atmosphere.given.file_option = "atmosphere_given_file";
    pism_config:atmosphere.given.file_type = "string";

    pism_config:atmosphere.given.periodic = "no";
    pism_config:atmosphere.given.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.given.periodic_type = "flag";

    pism_config:atmosphere.models = "given";
    pism_config:atmosphere.models_doc = "Comma-separated list of atmosphere melt models and modifiers";
    pism_config:atmosphere.models_option = "atmosphere";
    pism_config:atmosphere.models_type = "string";

    pism_config:atmosphere.one_station.file = "";
    pism_config:atmosphere.one_station.file_doc = "Specifies a file containing scalar time-series :var:`precipitation` and :var:`air_temp`.";
    pism_config:atmosphere.one_station.file_option = "atmosphere_one_station_file";
    pism_config:atmosphere.one_station.file_type = "string";

    pism_config:atmosphere.orographic_precipitation.background_precip_post = 0;
    pism_config:atmosphere.orographic_precipitation.background_precip_post_doc = "Background precipitation `P_{\\mathrm{post}}` added after the truncation.";
    pism_config:atmosphere.orographic_precipitation.background_precip_post_option = "background_precip_post";
    pism_config:atmosphere.orographic_precipitation.background_precip_post_type = "number";
    pism_config:atmosphere.orographic_precipitation.background_precip_post_units = "mm/hr";

    pism_config:atmosphere.orographic_precipitation.background_precip_pre = 0;
    pism_config:atmosphere.orographic_precipitation.background_precip_pre_doc = "Background precipitation `P_{\\mathrm{pre}}` added before the truncation.";
    pism_config:atmosphere.orographic_precipitation.background_precip_pre_option = "background_precip_pre";
    pism_config:atmosphere.orographic_precipitation.background_precip_pre_type = "number";
    pism_config:atmosphere.orographic_precipitation.background_precip_pre_units = "mm/hr";

    pism_config:atmosphere.orographic_precipitation.conversion_time = 1000.0;
    pism_config:atmosphere.orographic_precipitation.conversion_time_doc = "Cloud conversion time `\\tau_c`";
    pism_config:atmosphere.orographic_precipitation.conversion_time_option = "conversion_time";
    pism_config:atmosphere.orographic_precipitation.conversion_time_type = "number";
    pism_config:atmosphere.orographic_precipitation.conversion_time_units = "s";

    pism_config:atmosphere.orographic_precipitation.coriolis_latitude = 0.0;
    pism_config:atmosphere.orographic_precipitation.coriolis_latitude_doc = "Latitude used to compute Coriolis force";
    pism_config:atmosphere.orographic_precipitation.coriolis_latitude_option = "coriolis_latitude";
    pism_config:atmosphere.orographic_precipitation.coriolis_latitude_type = "number";
    pism_config:atmosphere.orographic_precipitation.coriolis_latitude_units = "degrees_N";

    pism_config:atmosphere.orographic_precipitation.fallout_time = 1000.0;
    pism_config:atmosphere.orographic_precipitation.fallout_time_doc = "Fallout time `\\tau_f`";
    pism_config:atmosphere.orographic_precipitation.fallout_time_option = "fallout_time";
    pism_config:atmosphere.orographic_precipitation.fallout_time_type = "number";
    pism_config:atmosphere.orographic_precipitation.fallout_time_units = "s";

    pism_config:atmosphere.orographic_precipitation.grid_size_factor = 2;
    pism_config:atmosphere.orographic_precipitation.grid_size_factor_doc = "The size of the extended grid is ``(Z*(grid.Mx - 1) + 1, Z*(grid.My - 1) + 1)`` where ``Z`` is given by this parameter.";
    pism_config:atmosphere.orographic_precipitation.grid_size_factor_type = "integer";
    pism_config:atmosphere.orographic_precipitation.grid_size_factor_units = "count";

    pism_config:atmosphere.orographic_precipitation.lapse_rate = -5.8;
    pism_config:atmosphere.orographic_precipitation.lapse_rate_doc = "Lapse rate `\\gamma`";
    pism_config:atmosphere.orographic_precipitation.lapse_rate_option = "lapse_rate";
    pism_config:atmosphere.orographic_precipitation.lapse_rate_type = "number";
    pism_config:atmosphere.orographic_precipitation.lapse_rate_units = "K / km";

    pism_config:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate = -6.5;
    pism_config:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_doc = "Moist adiabatic lapse rate `\\Gamma_m`";
    pism_config:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_option = "moist_adiabatic_lapse_rate";
    pism_config:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_type = "number";
    pism_config:atmosphere.orographic_precipitation.moist_adiabatic_lapse_rate_units = "K / km";

    pism_config:atmosphere.orographic_precipitation.moist_stability_frequency = 0.05;
    pism_config:atmosphere.orographic_precipitation.moist_stability_frequency_doc = "Moist stability frequency `N_m`";
    pism_config:atmosphere.orographic_precipitation.moist_stability_frequency_option = "moist_stability_frequency";
    pism_config:atmosphere.orographic_precipitation.moist_stability_frequency_type = "number";
    pism_config:atmosphere.orographic_precipitation.moist_stability_frequency_units = "1/s";

    pism_config:atmosphere.orographic_precipitation.reference_density = 7.4e-3;
    pism_config:atmosphere.orographic_precipitation.reference_density_doc = "Reference density `\\rho_{S_{\\text{ref}}}`";
    pism_config:atmosphere.orographic_precipitation.reference_density_option = "reference_density";
    pism_config:atmosphere.orographic_precipitation.reference_density_type = "number";
    pism_config:atmosphere.orographic_precipitation.reference_density_units = "kg m-3";

    pism_config:atmosphere.orographic_precipitation.scale_factor = 1;
    pism_config:atmosphere.orographic_precipitation.scale_factor_doc = "Precipitation scaling factor `S`.";
    pism_config:atmosphere.orographic_precipitation.scale_factor_option = "scale_factor";
    pism_config:atmosphere.orographic_precipitation.scale_factor_type = "number";
    pism_config:atmosphere.orographic_precipitation.scale_factor_units = "1";

    pism_config:atmosphere.orographic_precipitation.smoothing_standard_deviation = 0.0;
    pism_config:atmosphere.orographic_precipitation.smoothing_standard_deviation_doc = "Standard deviation of the Gaussian filter used to smooth surface elevation or zero if disabled";
    pism_config:atmosphere.orographic_precipitation.smoothing_standard_deviation_type = "number";
    pism_config:atmosphere.orographic_precipitation.smoothing_standard_deviation_units = "m";

    pism_config:atmosphere.orographic_precipitation.truncate = "true";
    pism_config:atmosphere.orographic_precipitation.truncate_doc = "Truncate precipitation at 0, disallowing negative precipitation values.";
    pism_config:atmosphere.orographic_precipitation.truncate_option = "truncate";
    pism_config:atmosphere.orographic_precipitation.truncate_type = "flag";

    pism_config:atmosphere.orographic_precipitation.water_vapor_scale_height = 2500.0;
    pism_config:atmosphere.orographic_precipitation.water_vapor_scale_height_doc = "Water vapor scale height `H_w`";
    pism_config:atmosphere.orographic_precipitation.water_vapor_scale_height_option = "water_vapor_scale_height";
    pism_config:atmosphere.orographic_precipitation.water_vapor_scale_height_type = "number";
    pism_config:atmosphere.orographic_precipitation.water_vapor_scale_height_units = "m";

    pism_config:atmosphere.orographic_precipitation.wind_direction = 270;
    pism_config:atmosphere.orographic_precipitation.wind_direction_doc = "The direction the wind is coming from";
    pism_config:atmosphere.orographic_precipitation.wind_direction_option = "wind_direction";
    pism_config:atmosphere.orographic_precipitation.wind_direction_type = "number";
    pism_config:atmosphere.orographic_precipitation.wind_direction_units = "degrees";

    pism_config:atmosphere.orographic_precipitation.wind_speed = 10;
    pism_config:atmosphere.orographic_precipitation.wind_speed_doc = "The wind speed.";
    pism_config:atmosphere.orographic_precipitation.wind_speed_option = "wind_speed";
    pism_config:atmosphere.orographic_precipitation.wind_speed_type = "number";
    pism_config:atmosphere.orographic_precipitation.wind_speed_units = "m/s";

    pism_config:atmosphere.pik.file = "";
    pism_config:atmosphere.pik.file_doc = "Name of the file containing the reference surface elevation field (variable :var:`usurf`).";
    pism_config:atmosphere.pik.file_option = "atmosphere_pik_file";
    pism_config:atmosphere.pik.file_type = "string";

    pism_config:atmosphere.pik.parameterization = "martin";
    pism_config:atmosphere.pik.parameterization_choices = "martin,huybrechts_dewolde,martin_huybrechts_dewolde,era_interim,era_interim_sin,era_interim_lon";
    pism_config:atmosphere.pik.parameterization_doc = "Selects parameterizations of mean annual and mean summer near-surface air temperatures.";
    pism_config:atmosphere.pik.parameterization_option = "atmosphere_pik";
    pism_config:atmosphere.pik.parameterization_type = "keyword";

    pism_config:atmosphere.precip_exponential_factor_for_temperature = 0.07041666667;
    pism_config:atmosphere.precip_exponential_factor_for_temperature_doc = "= 0.169/2.4; in SeaRISE-Greenland formula for precipitation correction using air temperature offsets relative to present; a 7.3\% change of precipitation rate for every one degC of temperature change :cite:`Huybrechts02`";
    pism_config:atmosphere.precip_exponential_factor_for_temperature_type = "number";
    pism_config:atmosphere.precip_exponential_factor_for_temperature_units = "Kelvin-1";

    pism_config:atmosphere.precip_scaling.file = "";
    pism_config:atmosphere.precip_scaling.file_doc = "Name of the file containing temperature offsets to use for a precipitation correction.";
    pism_config:atmosphere.precip_scaling.file_option = "atmosphere_precip_scaling_file";
    pism_config:atmosphere.precip_scaling.file_type = "string";

    pism_config:atmosphere.precip_scaling.periodic = "no";
    pism_config:atmosphere.precip_scaling.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.precip_scaling.periodic_type = "flag";

    pism_config:atmosphere.searise_greenland.file = "";
    pism_config:atmosphere.searise_greenland.file_doc = "Name of the file containing a precipitation field.";
    pism_config:atmosphere.searise_greenland.file_option = "atmosphere_searise_greenland_file";
    pism_config:atmosphere.searise_greenland.file_type = "string";

    pism_config:atmosphere.uniform.precipitation = 1000;
    pism_config:atmosphere.uniform.precipitation_doc = "Precipitation used by the ``uniform`` atmosphere model.";
    pism_config:atmosphere.uniform.precipitation_type = "number";
    pism_config:atmosphere.uniform.precipitation_units = "kg m-2 year-1";

    pism_config:atmosphere.uniform.temperature = 273.15;
    pism_config:atmosphere.uniform.temperature_doc = "Air temperature used by the ``uniform`` atmosphere model.";
    pism_config:atmosphere.uniform.temperature_type = "number";
    pism_config:atmosphere.uniform.temperature_units = "Kelvin";

    pism_config:atmosphere.yearly_cycle.file = "";
    pism_config:atmosphere.yearly_cycle.file_doc = "Name of the file containing mean annual and mean July temperatures (:var:`air_temp_mean_annual` and :var:`air_temp_mean_summer`) and the :var:`precipitation` field.";
    pism_config:atmosphere.yearly_cycle.file_option = "atmosphere_yearly_cycle_file";
    pism_config:atmosphere.yearly_cycle.file_type = "string";

    pism_config:atmosphere.yearly_cycle.scaling.file = "";
    pism_config:atmosphere.yearly_cycle.scaling.file_doc = "Name of the file containing amplitude scaling (:var:`amplitude_scaling`) for the near-surface air temperature.";
    pism_config:atmosphere.yearly_cycle.scaling.file_option = "atmosphere_yearly_cycle_scaling_file";
    pism_config:atmosphere.yearly_cycle.scaling.file_type = "string";

    pism_config:atmosphere.yearly_cycle.scaling.periodic = "no";
    pism_config:atmosphere.yearly_cycle.scaling.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:atmosphere.yearly_cycle.scaling.periodic_type = "flag";

    pism_config:basal_resistance.beta_ice_free_bedrock = 1.8e9;
    pism_config:basal_resistance.beta_ice_free_bedrock_doc = "value is for ice stream E from :cite:`HulbeMacAyeal`; thus sliding velocity, but we hope it doesn't matter much; at 100 m/year the linear sliding law gives 57040 Pa basal shear stress";
    pism_config:basal_resistance.beta_ice_free_bedrock_type = "number";
    pism_config:basal_resistance.beta_ice_free_bedrock_units = "Pascal second meter-1";

    pism_config:basal_resistance.beta_lateral_margin = 1e19;
    pism_config:basal_resistance.beta_lateral_margin_doc = "high value of `\\beta` used to simulate drag at lateral ice margins (fjord walls, etc); the default value is chosen to disable flow in the direction along a margin";
    pism_config:basal_resistance.beta_lateral_margin_type = "number";
    pism_config:basal_resistance.beta_lateral_margin_units = "Pascal second meter-1";

    pism_config:basal_resistance.plastic.regularization = 0.01;
    pism_config:basal_resistance.plastic.regularization_doc = "Set the value of `\\epsilon` regularization of plastic till; this is the second `\\epsilon` in formula (4.1) in :cite:`SchoofStream`";
    pism_config:basal_resistance.plastic.regularization_option = "plastic_reg";
    pism_config:basal_resistance.plastic.regularization_type = "number";
    pism_config:basal_resistance.plastic.regularization_units = "meter / year";

    pism_config:basal_resistance.pseudo_plastic.enabled = "no";
    pism_config:basal_resistance.pseudo_plastic.enabled_doc = "Use the pseudo-plastic till model (basal sliding law).";
    pism_config:basal_resistance.pseudo_plastic.enabled_option = "pseudo_plastic";
    pism_config:basal_resistance.pseudo_plastic.enabled_type = "flag";

    pism_config:basal_resistance.pseudo_plastic.q = 0.25;
    pism_config:basal_resistance.pseudo_plastic.q_doc = "The exponent of the pseudo-plastic basal resistance model";
    pism_config:basal_resistance.pseudo_plastic.q_option = "pseudo_plastic_q";
    pism_config:basal_resistance.pseudo_plastic.q_type = "number";
    pism_config:basal_resistance.pseudo_plastic.q_units = "pure number";

    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor = -1.0;
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_doc = "divides pseudo-plastic tauc (yield stress) by given factor; this would increase sliding by given factor in absence of membrane stresses; not used if negative or zero; not used by default";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_option = "sliding_scale_factor_reduces_tauc";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_type = "number";
    pism_config:basal_resistance.pseudo_plastic.sliding_scale_factor_units = "1";

    pism_config:basal_resistance.pseudo_plastic.u_threshold = 100.0;
    pism_config:basal_resistance.pseudo_plastic.u_threshold_doc = "threshold velocity of the pseudo-plastic sliding law";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_option = "pseudo_plastic_uthreshold";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_type = "number";
    pism_config:basal_resistance.pseudo_plastic.u_threshold_units = "meter / year";

    pism_config:basal_resistance.regularized_coulomb.enabled = "no";
    pism_config:basal_resistance.regularized_coulomb.enabled_doc = "Use the regularized Coulomb till friction model (basal sliding law) as in equation (3) in :cite:`ZoetIverson20`";
    pism_config:basal_resistance.regularized_coulomb.enabled_option = "regularized_coulomb";
    pism_config:basal_resistance.regularized_coulomb.enabled_type = "flag";

    pism_config:basal_yield_stress.add_transportable_water = "no";
    pism_config:basal_yield_stress.add_transportable_water_doc = "If \"yes\" then the water amount in the transport system is added to tillwat in determining tauc (in the Mohr-Coulomb relation).  Normally only the water in the till is used.";
    pism_config:basal_yield_stress.add_transportable_water_option = "tauc_add_transportable_water";
    pism_config:basal_yield_stress.add_transportable_water_type = "flag";

    pism_config:basal_yield_stress.constant.value = 2e5;
    pism_config:basal_yield_stress.constant.value_doc = "fill value for yield stress for basal till (plastic or pseudo-plastic model); note `2 \\times 10^5` Pa = 2 bar is quite strong and little sliding should occur";
    pism_config:basal_yield_stress.constant.value_option = "tauc";
    pism_config:basal_yield_stress.constant.value_type = "number";
    pism_config:basal_yield_stress.constant.value_units = "Pascal";

    pism_config:basal_yield_stress.ice_free_bedrock = 1e6;
    pism_config:basal_yield_stress.ice_free_bedrock_doc = "the \"high\" yield stress value used in grounded ice-free areas.";
    pism_config:basal_yield_stress.ice_free_bedrock_option = "high_tauc";
    pism_config:basal_yield_stress.ice_free_bedrock_type = "number";
    pism_config:basal_yield_stress.ice_free_bedrock_units = "Pascal";

    pism_config:basal_yield_stress.model = "mohr_coulomb";
    pism_config:basal_yield_stress.model_choices = "constant,mohr_coulomb,tillphi_opt";
    pism_config:basal_yield_stress.model_doc = "The basal yield stress model to use when sliding is active.";
    pism_config:basal_yield_stress.model_option = "yield_stress";
    pism_config:basal_yield_stress.model_type = "keyword";

    pism_config:basal_yield_stress.mohr_coulomb.delta.file = "";
    pism_config:basal_yield_stress.mohr_coulomb.delta.file_doc = "Name of the file containing space- and time-dependent variable :var:`mohr_coulomb_delta` to use instead of :config:`basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden`.";
    pism_config:basal_yield_stress.mohr_coulomb.delta.file_option = "mohr_coulomb_delta_file";
    pism_config:basal_yield_stress.mohr_coulomb.delta.file_type = "string";

    pism_config:basal_yield_stress.mohr_coulomb.delta.periodic = "no";
    pism_config:basal_yield_stress.mohr_coulomb.delta.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:basal_yield_stress.mohr_coulomb.delta.periodic_type = "flag";

    pism_config:basal_yield_stress.mohr_coulomb.tauc_to_phi.file = "";
    pism_config:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_doc = "File containing the basal yield stress field that should be used to recover the till friction angle distribution.";
    pism_config:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_option = "tauc_to_phi";
    pism_config:basal_yield_stress.mohr_coulomb.tauc_to_phi.file_type = "string";

    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion = 0.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_doc = "cohesion of till; = `c_0` in most references; note Schoof uses zero but Paterson pp 168--169 gives range 0--40 kPa; but Paterson notes that \"... all the pairs `c_0` and `\\phi` in the table would give a yield stress for Ice Stream B that exceeds the basal shear stress there...\"";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_option = "till_cohesion";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_cohesion_units = "Pascal";

    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient = 0.12;
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_doc = "coefficient of compressiblity of till; value from :cite:`Tulaczyketal2000`";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_option = "till_compressibility_coefficient";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_compressibility_coefficient_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden = 0.02;
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_doc = "`\\delta` in :cite:`BuelervanPelt2015`; `\\delta P_o \\le N_{\\text{till}} \\le P_o` where `P_o` is overburden pressure and `N_{\\text{till}}` is the effective pressure of the overlying ice on the saturated till; default value of `\\delta` corresponds to  Greenland and Antarctic model runs";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_option = "till_effective_fraction_overburden";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water = 0.1;
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_doc = "If :config:`basal_yield_stress.add_transportable_water` is set then the water amount in the transport system is added to :var:`tillwat` in determining :var:`tauc`.  Normally only the water in the till is used.  This factor multiplies the logarithm in that formula.";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_option = "till_log_factor_transportable_water";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_log_factor_transportable_water_units = "meters";

    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default = 30.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_doc = "fill value for till friction angle";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_option = "plastic_phi";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_phi_default_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure = 1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_doc = "reference effective pressure `N_0`; value from :cite:`Tulaczyketal2000`";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_effective_pressure_units = "Pascal";

    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio = 0.69;
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_doc = "void ratio at reference effective pressure `N_0`; value from :cite:`Tulaczyketal2000`";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_option = "till_reference_void_ratio";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.till_reference_void_ratio_units = "pure number";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dhdt_min = 0.001;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dhdt_min_doc = "rate of change in the surface elevation mismatch `D` used as a convergence criterion";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dhdt_min_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dhdt_min_units = "meters year-1";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dhdt_min_option = "tillphi_opt_dhdt_min";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_max = 1.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_max_doc = "maximum till friction angle adjustment `\\dphimax`";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_max_units = "degrees";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_max_option = "tillphi_opt_dphi_max";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_scale = 2e-3;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_scale_doc = "scaling factor `C` used to compute the `\\Delta \\phi` adjustment, `C` degrees per meter of surface elevation mismatch";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_scale_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_scale_units = "degree / meters";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dphi_scale_option = "tillphi_opt_dphi_scale";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dt = 250.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dt_doc = "time step `\\dt_{\\phi}` for optimization of till friction angle";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dt_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dt_units = "365days";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.dt_option = "tillphi_opt_dt";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.file = "";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.file_doc = "Name of the file containing the time-independent variable :var:`usurf` used as target surface elevation";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.file_option = "tillphi_opt_file";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.file_type = "string";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max = 5.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max_doc = "maximum value of the lower bound of the till friction angle, `\\phi_{0,\\mathrm{max}}`";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max_units = "degrees";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max_option = "tillphi_opt_phi0_max";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min = 2.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min_doc = "minimum value of the lower bound of the till friction angle, `\\phi_{0,\\mathrm{min}}`";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min_units = "degrees";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min_option = "tillphi_opt_phi0_min";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi_max = 70.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi_max_doc = "upper bound of the till friction angle `\\phimax`";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi_max_units = "degrees";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.phi_max_option = "tillphi_opt_phi_max";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_max = 700.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_max_doc = "the bed elevation `\\bmax` above which :config:`basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_max` is used";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_max_units = "meters";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_max_option = "tillphi_opt_topg_max";

    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_min = -300.0;
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_min_doc = "the bed elevation `\\bmin` below which :config:`basal_yield_stress.mohr_coulomb.tillphi_opt.phi0_min` is used";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_min_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_min_units = "meters";
    pism_config:basal_yield_stress.mohr_coulomb.tillphi_opt.topg_min_option = "tillphi_opt_topg_min";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled = "no";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_doc = "If the option ``-topg_to_phi`` is set then this will be set to \"yes\", and then ``MohrCoulombYieldStress`` will initialize the :var:`tillphi` field using a piece-wise linear function of depth described by four parameters.";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled_type = "flag";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max = 15.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_doc = "upper value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min = 5.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_doc = "lower value of the till friction angle; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min_units = "degrees";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max = 1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_doc = "the elevation at which the upper value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max_units = "meters";

    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min = -1000.0;
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_doc = "the elevation at which the lower value of the till friction angle is used; see the implementation of MohrCoulombYieldStress";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_type = "number";
    pism_config:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min_units = "meters";

    pism_config:basal_yield_stress.slippery_grounding_lines = "no";
    pism_config:basal_yield_stress.slippery_grounding_lines_doc = "If yes, at icy grounded locations with bed elevations below sea level, within one cell of floating ice or ice-free ocean, make tauc as low as possible from the Mohr-Coulomb relation.  Specifically, at such locations replace the normally-computed tauc from the Mohr-Coulomb relation, which uses the effective pressure from the modeled amount of water in the till, by the minimum value of tauc from Mohr-Coulomb, i.e. by using the effective pressure corresponding to the maximum amount of till-stored water.  Does not alter the modeled or reported amount of till water, nor does this mechanism affect water conservation.";
    pism_config:basal_yield_stress.slippery_grounding_lines_option = "tauc_slippery_grounding_lines";
    pism_config:basal_yield_stress.slippery_grounding_lines_type = "flag";

    pism_config:bed_deformation.bed_topography_delta_file = "";
    pism_config:bed_deformation.bed_topography_delta_file_doc = "The name of the file to read the :var:`topg_delta` from. This field is added to the bed topography during initialization.";
    pism_config:bed_deformation.bed_topography_delta_file_option = "topg_delta_file";
    pism_config:bed_deformation.bed_topography_delta_file_type = "string";

    pism_config:bed_deformation.bed_uplift_file = "";
    pism_config:bed_deformation.bed_uplift_file_doc = "The name of the file to read the uplift (dbdt) from. Leave empty to read it from an input file or a regridding file.";
    pism_config:bed_deformation.bed_uplift_file_option = "uplift_file";
    pism_config:bed_deformation.bed_uplift_file_type = "string";

    pism_config:bed_deformation.given.file = "";
    pism_config:bed_deformation.given.file_doc = "Name of the file containing time-dependent :var:`topg_delta`.";
    pism_config:bed_deformation.given.file_option = "topg_delta_file";
    pism_config:bed_deformation.given.file_type = "string";

    pism_config:bed_deformation.given.reference_file = "";
    pism_config:bed_deformation.given.reference_file_doc = "Name of the file containing the reference bed topography :var:`topg`.";
    pism_config:bed_deformation.given.reference_file_option = "topg_reference_file";
    pism_config:bed_deformation.given.reference_file_type = "string";

    pism_config:bed_deformation.lc.elastic_model = "yes";
    pism_config:bed_deformation.lc.elastic_model_doc = "Use the elastic part of the Lingle-Clark bed deformation model.";
    pism_config:bed_deformation.lc.elastic_model_option = "bed_def_lc_elastic_model";
    pism_config:bed_deformation.lc.elastic_model_type = "flag";

    pism_config:bed_deformation.lc.grid_size_factor = 4;
    pism_config:bed_deformation.lc.grid_size_factor_doc = "The spectral grid size is ``(Z*(grid.Mx - 1) + 1, Z*(grid.My - 1) + 1)`` where ``Z`` is given by this parameter. See :cite:`LingleClark`, :cite:`BLKfastearth`.";
    pism_config:bed_deformation.lc.grid_size_factor_type = "integer";
    pism_config:bed_deformation.lc.grid_size_factor_units = "count";

    pism_config:bed_deformation.lc.update_interval = 10.0;
    pism_config:bed_deformation.lc.update_interval_doc = "Interval between updates of the Lingle-Clark model";
    pism_config:bed_deformation.lc.update_interval_type = "number";
    pism_config:bed_deformation.lc.update_interval_units = "365days";

    pism_config:bed_deformation.lithosphere_flexural_rigidity = 5.0e24;
    pism_config:bed_deformation.lithosphere_flexural_rigidity_doc = "lithosphere flexural rigidity used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_config:bed_deformation.lithosphere_flexural_rigidity_type = "number";
    pism_config:bed_deformation.lithosphere_flexural_rigidity_units = "Newton meter";

    pism_config:bed_deformation.mantle_density = 3300.0;
    pism_config:bed_deformation.mantle_density_doc = "half-space (mantle) density used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_config:bed_deformation.mantle_density_type = "number";
    pism_config:bed_deformation.mantle_density_units = "kg meter-3";

    pism_config:bed_deformation.mantle_viscosity = 1.0e21;
    pism_config:bed_deformation.mantle_viscosity_doc = "half-space (mantle) viscosity used by the bed deformation model. See :cite:`LingleClark`, :cite:`BLKfastearth`";
    pism_config:bed_deformation.mantle_viscosity_type = "number";
    pism_config:bed_deformation.mantle_viscosity_units = "Pascal second";

    pism_config:bed_deformation.model = "none";
    pism_config:bed_deformation.model_choices = "none,iso,lc,given";
    pism_config:bed_deformation.model_doc = "Selects a bed deformation model to use. ``iso`` is point-wise isostasy, ``lc`` is the Lingle-Clark model (see :cite:`LingleClark`, requires FFTW_), ``given`` uses prescribed bed topography changes read from a file.";
    pism_config:bed_deformation.model_option = "bed_def";
    pism_config:bed_deformation.model_type = "keyword";

    pism_config:bootstrapping.defaults.bed = 1.0;
    pism_config:bootstrapping.defaults.bed_doc = "bed elevation value to use if :var:`topg` (``bedrock_altitude``) variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bed_type = "number";
    pism_config:bootstrapping.defaults.bed_units = "meters";

    pism_config:bootstrapping.defaults.bmelt = 0.0;
    pism_config:bootstrapping.defaults.bmelt_doc = "basal melt rate value to use if variable :var:`bmelt` is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bmelt_type = "number";
    pism_config:bootstrapping.defaults.bmelt_units = "meter / second";

    pism_config:bootstrapping.defaults.bwat = 0.0;
    pism_config:bootstrapping.defaults.bwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.bwat_type = "number";
    pism_config:bootstrapping.defaults.bwat_units = "meters";

    pism_config:bootstrapping.defaults.bwp = 0.0;
    pism_config:bootstrapping.defaults.bwp_doc = "basal water pressure value to use if variable :var:`bwp` is absent in bootstrapping file; most hydrology models do not use this value because :var:`bwp` is diagnostic";
    pism_config:bootstrapping.defaults.bwp_type = "number";
    pism_config:bootstrapping.defaults.bwp_units = "Pascal";

    pism_config:bootstrapping.defaults.geothermal_flux = 0.042;
    pism_config:bootstrapping.defaults.geothermal_flux_doc = "geothermal flux value to use if bheatflx variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.geothermal_flux_type = "number";
    pism_config:bootstrapping.defaults.geothermal_flux_units = "Watt meter-2";

    pism_config:bootstrapping.defaults.ice_thickness = 0.0;
    pism_config:bootstrapping.defaults.ice_thickness_doc = "thickness value to use if thk (land_ice_thickness) variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.ice_thickness_type = "number";
    pism_config:bootstrapping.defaults.ice_thickness_units = "meters";

    pism_config:bootstrapping.defaults.tillwat = 0.0;
    pism_config:bootstrapping.defaults.tillwat_doc = "till water thickness value to use if variable tillwat is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.tillwat_type = "number";
    pism_config:bootstrapping.defaults.tillwat_units = "meters";

    pism_config:bootstrapping.defaults.uplift = 0.0;
    pism_config:bootstrapping.defaults.uplift_doc = "uplift value to use if dbdt variable is absent in bootstrapping file";
    pism_config:bootstrapping.defaults.uplift_type = "number";
    pism_config:bootstrapping.defaults.uplift_units = "meter / second";

    pism_config:bootstrapping.temperature_heuristic = "smb";
    pism_config:bootstrapping.temperature_heuristic_choices = "smb,quartic_guess";
    pism_config:bootstrapping.temperature_heuristic_doc = "The heuristic to use to initialize ice temperature during bootstrapping: ``smb`` uses the surface mass balance, surface temperature, and the geothermal flux, ``quartic_guess`` uses the surface temperature and the geothermal flux.";
    pism_config:bootstrapping.temperature_heuristic_option = "boot_temperature_heuristic";
    pism_config:bootstrapping.temperature_heuristic_type = "keyword";

    pism_config:calving.eigen_calving.K = 0.0;
    pism_config:calving.eigen_calving.K_doc = "Set proportionality constant to determine calving rate from strain rates.  Note references :cite:`Levermannetal2012`, :cite:`Martinetal2011` use K in range `10^{9}` to `3 \\times 10^{11}` m a, that is, `3 \\times 10^{16}` to `10^{19}` m s.";
    pism_config:calving.eigen_calving.K_option = "eigen_calving_K";
    pism_config:calving.eigen_calving.K_type = "number";
    pism_config:calving.eigen_calving.K_units = "meter second";

    pism_config:calving.float_kill.calve_near_grounding_line = "yes";
    pism_config:calving.float_kill.calve_near_grounding_line_doc = "Calve floating ice near the grounding line.";
    pism_config:calving.float_kill.calve_near_grounding_line_option = "float_kill_calve_near_grounding_line";
    pism_config:calving.float_kill.calve_near_grounding_line_type = "flag";

    pism_config:calving.float_kill.margin_only = "no";
    pism_config:calving.float_kill.margin_only_doc = "Apply float_kill at ice margin cells only.";
    pism_config:calving.float_kill.margin_only_option = "float_kill_margin_only";
    pism_config:calving.float_kill.margin_only_type = "flag";

    pism_config:calving.hayhurst_calving.B_tilde = 65.0;
    pism_config:calving.hayhurst_calving.B_tilde_doc = "Effective damage rate :cite:`Mercenier2018`";
    pism_config:calving.hayhurst_calving.B_tilde_type = "number";
    pism_config:calving.hayhurst_calving.B_tilde_units = "(MPa)^r / year";

    pism_config:calving.hayhurst_calving.exponent_r = 0.43;
    pism_config:calving.hayhurst_calving.exponent_r_doc = "Damage law exponent :cite:`Mercenier2018`";
    pism_config:calving.hayhurst_calving.exponent_r_type = "number";
    pism_config:calving.hayhurst_calving.exponent_r_units = "1";

    pism_config:calving.hayhurst_calving.sigma_threshold = 0.17;
    pism_config:calving.hayhurst_calving.sigma_threshold_doc = "Damage threshold stress :cite:`Mercenier2018`";
    pism_config:calving.hayhurst_calving.sigma_threshold_type = "number";
    pism_config:calving.hayhurst_calving.sigma_threshold_units = "MPa";

    pism_config:calving.methods = "";
    pism_config:calving.methods_doc = "comma-separated list of calving methods; one or more of ``eigen_calving``, ``float_kill``, ``thickness_calving``";
    pism_config:calving.methods_option = "calving";
    pism_config:calving.methods_type = "string";

    pism_config:calving.rate_scaling.file = "";
    pism_config:calving.rate_scaling.file_doc = "File containing the scaling factor applied to calving rates from ``eigen_calving``, ``vonmises_calving``, and ``hayhurst_calving`` (variable name: ``frac_calving_rate``)";
    pism_config:calving.rate_scaling.file_type = "string";

    pism_config:calving.rate_scaling.periodic = "no";
    pism_config:calving.rate_scaling.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:calving.rate_scaling.periodic_type = "flag";

    pism_config:calving.thickness_calving.file = "";
    pism_config:calving.thickness_calving.file_doc = "Name of the file containing the spatially-variable thickness calving threshold.";
    pism_config:calving.thickness_calving.file_option = "thickness_calving_file";
    pism_config:calving.thickness_calving.file_type = "string";

    pism_config:calving.thickness_calving.periodic = "no";
    pism_config:calving.thickness_calving.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:calving.thickness_calving.periodic_type = "flag";

    pism_config:calving.thickness_calving.threshold = 50.0;
    pism_config:calving.thickness_calving.threshold_doc = "When terminal ice thickness of floating ice shelf is less than this threshold, it will be calved off.";
    pism_config:calving.thickness_calving.threshold_option = "thickness_calving_threshold";
    pism_config:calving.thickness_calving.threshold_type = "number";
    pism_config:calving.thickness_calving.threshold_units = "meters";

    pism_config:calving.vonmises_calving.Glen_exponent = 3.0;
    pism_config:calving.vonmises_calving.Glen_exponent_doc = "Glen exponent in ice flow law for von Mises calving";
    pism_config:calving.vonmises_calving.Glen_exponent_option = "vonmises_calving_n";
    pism_config:calving.vonmises_calving.Glen_exponent_type = "number";
    pism_config:calving.vonmises_calving.Glen_exponent_units = "pure number";

    pism_config:calving.vonmises_calving.flow_law = "gpbld";
    pism_config:calving.vonmises_calving.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb";
    pism_config:calving.vonmises_calving.flow_law_doc = "The custom flow law for the von Mises stress computation";
    pism_config:calving.vonmises_calving.flow_law_type = "keyword";

    pism_config:calving.vonmises_calving.sigma_max = 1.0e6;
    pism_config:calving.vonmises_calving.sigma_max_doc = "Set maximum tensile stress.  Note references :cite:`Morlighem2016` use 1.0e6 Pa.";
    pism_config:calving.vonmises_calving.sigma_max_option = "vonmises_calving_calving_sigma_max";
    pism_config:calving.vonmises_calving.sigma_max_type = "number";
    pism_config:calving.vonmises_calving.sigma_max_units = "Pa";

    pism_config:calving.vonmises_calving.threshold_file = "";
    pism_config:calving.vonmises_calving.threshold_file_doc = "Name of the file containing the spatially-variable :var:`vonmises_calving_threshold`.";
    pism_config:calving.vonmises_calving.threshold_file_option = "vonmises_calving_threshold_file";
    pism_config:calving.vonmises_calving.threshold_file_type = "string";

    pism_config:calving.vonmises_calving.use_custom_flow_law = "no";
    pism_config:calving.vonmises_calving.use_custom_flow_law_doc = "Use custom flow law in the von Mises stress computation";
    pism_config:calving.vonmises_calving.use_custom_flow_law_option = "vonmises_calving_use_custom_flow_law";
    pism_config:calving.vonmises_calving.use_custom_flow_law_type = "flag";

    pism_config:constants.fresh_water.density = 1000.0;
    pism_config:constants.fresh_water.density_doc = "density of fresh water";
    pism_config:constants.fresh_water.density_type = "number";
    pism_config:constants.fresh_water.density_units = "kg meter-3";

    pism_config:constants.fresh_water.latent_heat_of_fusion = 3.34e5;
    pism_config:constants.fresh_water.latent_heat_of_fusion_doc = "latent heat of fusion for water :cite:`AschwandenBlatter`";
    pism_config:constants.fresh_water.latent_heat_of_fusion_type = "number";
    pism_config:constants.fresh_water.latent_heat_of_fusion_units = "Joule / kg";

    pism_config:constants.fresh_water.melting_point_temperature = 273.15;
    pism_config:constants.fresh_water.melting_point_temperature_doc = "melting point of pure water";
    pism_config:constants.fresh_water.melting_point_temperature_type = "number";
    pism_config:constants.fresh_water.melting_point_temperature_units = "Kelvin";

    pism_config:constants.fresh_water.specific_heat_capacity = 4170.0;
    pism_config:constants.fresh_water.specific_heat_capacity_doc = "at melting point T_0 :cite:`AschwandenBlatter`";
    pism_config:constants.fresh_water.specific_heat_capacity_type = "number";
    pism_config:constants.fresh_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.global_ocean_area = 3.625e14;
    pism_config:constants.global_ocean_area_doc = "area of the global ocean :cite:`Cogley2011`";
    pism_config:constants.global_ocean_area_type = "number";
    pism_config:constants.global_ocean_area_units = "meter2";

    pism_config:constants.ice.beta_Clausius_Clapeyron = 7.9e-8;
    pism_config:constants.ice.beta_Clausius_Clapeyron_doc = "Clausius-Clapeyron constant relating melting temperature and pressure: `\\beta = dT / dP` :cite:`Luethi2002`";
    pism_config:constants.ice.beta_Clausius_Clapeyron_type = "number";
    pism_config:constants.ice.beta_Clausius_Clapeyron_units = "Kelvin / Pascal";

    pism_config:constants.ice.density = 910.0;
    pism_config:constants.ice.density_doc = "`\\rho_i`; density of ice in ice sheet";
    pism_config:constants.ice.density_type = "number";
    pism_config:constants.ice.density_units = "kg meter-3";

    pism_config:constants.ice.grain_size = 1.0;
    pism_config:constants.ice.grain_size_doc = "Default constant ice grain size to use with the Goldsby-Kohlstedt :cite:`GoldsbyKohlstedt` flow law";
    pism_config:constants.ice.grain_size_option = "ice_grain_size";
    pism_config:constants.ice.grain_size_type = "number";
    pism_config:constants.ice.grain_size_units = "mm";

    pism_config:constants.ice.specific_heat_capacity = 2009.0;
    pism_config:constants.ice.specific_heat_capacity_doc = "specific heat capacity of pure ice at melting point T_0";
    pism_config:constants.ice.specific_heat_capacity_type = "number";
    pism_config:constants.ice.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.ice.thermal_conductivity = 2.10;
    pism_config:constants.ice.thermal_conductivity_doc = "= W m-1 K-1; thermal conductivity of pure ice";
    pism_config:constants.ice.thermal_conductivity_type = "number";
    pism_config:constants.ice.thermal_conductivity_units = "Joule / (meter Kelvin second)";

    pism_config:constants.ideal_gas_constant = 8.31441;
    pism_config:constants.ideal_gas_constant_doc = "ideal gas constant";
    pism_config:constants.ideal_gas_constant_type = "number";
    pism_config:constants.ideal_gas_constant_units = "Joule / (mol Kelvin)";

    pism_config:constants.sea_water.density = 1028.0;
    pism_config:constants.sea_water.density_doc = "density of sea water";
    pism_config:constants.sea_water.density_type = "number";
    pism_config:constants.sea_water.density_units = "kg meter-3";

    pism_config:constants.sea_water.salinity = 35.0;
    pism_config:constants.sea_water.salinity_doc = "salinity of sea water";
    pism_config:constants.sea_water.salinity_type = "number";
    pism_config:constants.sea_water.salinity_units = "g / kg";

    pism_config:constants.sea_water.specific_heat_capacity = 3985.0;
    pism_config:constants.sea_water.specific_heat_capacity_doc = "at 35 psu, value taken from `Kaye and Laby`_, section 2.7.9";
    pism_config:constants.sea_water.specific_heat_capacity_type = "number";
    pism_config:constants.sea_water.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:constants.standard_gravity = 9.81;
    pism_config:constants.standard_gravity_doc = "acceleration due to gravity on Earth geoid";
    pism_config:constants.standard_gravity_type = "number";
    pism_config:constants.standard_gravity_units = "meter second-2";

    pism_config:energy.allow_temperature_above_melting = "no";
    pism_config:energy.allow_temperature_above_melting_doc = "If set to \"yes\", allow temperatures above the pressure-malting point in the cold mode temperature code. Used by some verifiaction tests.";
    pism_config:energy.allow_temperature_above_melting_type = "flag";

    pism_config:energy.basal_melt.use_grounded_cell_fraction  = "true";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_doc = "If geometry.grounded_cell_fraction is set, use the fractional floatation mask to interpolate the basal melt rate at the grounding line between grounded and floating values.";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_option  = "subgl_basal_melt";
    pism_config:energy.basal_melt.use_grounded_cell_fraction_type  = "flag";

    pism_config:energy.bedrock_thermal.conductivity = 3.0;
    pism_config:energy.bedrock_thermal.conductivity_doc = "= W m-1 K-1; for bedrock used in thermal model :cite:`RitzEISMINT`";
    pism_config:energy.bedrock_thermal.conductivity_type = "number";
    pism_config:energy.bedrock_thermal.conductivity_units = "Joule / (meter Kelvin second)";

    pism_config:energy.bedrock_thermal.density = 3300.0;
    pism_config:energy.bedrock_thermal.density_doc = "for bedrock used in thermal model";
    pism_config:energy.bedrock_thermal.density_type = "number";
    pism_config:energy.bedrock_thermal.density_units = "kg meter-3";

    pism_config:energy.bedrock_thermal.file = "";
    pism_config:energy.bedrock_thermal.file_doc = "Name of the file containing the geothermal flux field :var:`bheatflx`. Leave empty to read it from the :config:`input.file`.";
    pism_config:energy.bedrock_thermal.file_type = "string";

    pism_config:energy.bedrock_thermal.specific_heat_capacity = 1000.0;
    pism_config:energy.bedrock_thermal.specific_heat_capacity_doc = "for bedrock used in thermal model :cite:`RitzEISMINT`";
    pism_config:energy.bedrock_thermal.specific_heat_capacity_type = "number";
    pism_config:energy.bedrock_thermal.specific_heat_capacity_units = "Joule / (kg Kelvin)";

    pism_config:energy.ch_warming.average_channel_spacing = 20.0;
    pism_config:energy.ch_warming.average_channel_spacing_doc = "Average spacing between elements of the cryo-hydrologic system (controls the rate of heat transfer from the CH system into the ice).";
    pism_config:energy.ch_warming.average_channel_spacing_type = "number";
    pism_config:energy.ch_warming.average_channel_spacing_units = "meters";

    pism_config:energy.ch_warming.enabled = "no";
    pism_config:energy.ch_warming.enabled_doc = "Enable the cryo-hydrologic warming model";
    pism_config:energy.ch_warming.enabled_type = "flag";

    pism_config:energy.ch_warming.residual_water_fraction = 0.005;
    pism_config:energy.ch_warming.residual_water_fraction_doc = "residual water fraction in the cryo-hydrologic system at the end of a melt season";
    pism_config:energy.ch_warming.residual_water_fraction_type = "number";
    pism_config:energy.ch_warming.residual_water_fraction_units = "pure number";

    pism_config:energy.ch_warming.temperate_ice_thermal_conductivity_ratio = 1.0;
    pism_config:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_doc = "ratio of thermal conductivities of temperate and cold ice in the cryo-hydrologic system";
    pism_config:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_type = "number";
    pism_config:energy.ch_warming.temperate_ice_thermal_conductivity_ratio_units = "pure number";

    pism_config:energy.drainage_maximum_rate = 1.58443823077064e-09;
    pism_config:energy.drainage_maximum_rate_doc = "0.05 year-1; maximum rate at which liquid water fraction in temperate ice could possibly drain; see :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_config:energy.drainage_maximum_rate_type = "number";
    pism_config:energy.drainage_maximum_rate_units = "second-1";

    pism_config:energy.drainage_target_water_fraction = 0.01;
    pism_config:energy.drainage_target_water_fraction_doc = "liquid water fraction (omega) above which drainage occurs, but below which there is no drainage; see :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_config:energy.drainage_target_water_fraction_type = "number";
    pism_config:energy.drainage_target_water_fraction_units = "1";

    pism_config:energy.enabled = "yes";
    pism_config:energy.enabled_doc = "Solve energy conservation equations.";
    pism_config:energy.enabled_type = "flag";

    pism_config:energy.enthalpy.cold_bulge_max = 60270.0;
    pism_config:energy.enthalpy.cold_bulge_max_doc = "= (2009 J kg-1 K-1) * (30 K); maximum amount by which advection can reduce the enthalpy of a column of ice below its surface enthalpy value";
    pism_config:energy.enthalpy.cold_bulge_max_type = "number";
    pism_config:energy.enthalpy.cold_bulge_max_units = "Joule / kg";

    pism_config:energy.enthalpy.temperate_ice_thermal_conductivity_ratio = 0.1;
    pism_config:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_doc = "K in cold ice is multiplied by this fraction to give K0 in :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_config:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_type = "number";
    pism_config:energy.enthalpy.temperate_ice_thermal_conductivity_ratio_units = "pure number";

    pism_config:energy.margin_exclude_horizontal_advection = "yes";
    pism_config:energy.margin_exclude_horizontal_advection_doc = "Exclude horizontal advection of energy at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_config:energy.margin_exclude_horizontal_advection_type = "flag";

    pism_config:energy.margin_exclude_strain_heating = "yes";
    pism_config:energy.margin_exclude_strain_heating_doc = "Exclude strain heating at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_config:energy.margin_exclude_strain_heating_type = "flag";

    pism_config:energy.margin_exclude_vertical_advection = "yes";
    pism_config:energy.margin_exclude_vertical_advection_doc = "Exclude vertical advection of energy at grid points near ice margins. See :config:`energy.margin_ice_thickness_limit`.";
    pism_config:energy.margin_exclude_vertical_advection_type = "flag";

    pism_config:energy.margin_ice_thickness_limit = 100.0;
    pism_config:energy.margin_ice_thickness_limit_doc = "use special margin treatment at grid points with a neighbor with the thickness below this limit.";
    pism_config:energy.margin_ice_thickness_limit_type = "number";
    pism_config:energy.margin_ice_thickness_limit_units = "meters";

    pism_config:energy.max_low_temperature_count = 10;
    pism_config:energy.max_low_temperature_count_doc = "Maximum number of grid points with ice temperature below energy.minimum_allowed_temperature.";
    pism_config:energy.max_low_temperature_count_option = "max_low_temps";
    pism_config:energy.max_low_temperature_count_type = "integer";
    pism_config:energy.max_low_temperature_count_units = "count";

    pism_config:energy.minimum_allowed_temperature = 200.0;
    pism_config:energy.minimum_allowed_temperature_doc = "Minimum allowed ice temperature";
    pism_config:energy.minimum_allowed_temperature_option = "low_temp";
    pism_config:energy.minimum_allowed_temperature_type = "number";
    pism_config:energy.minimum_allowed_temperature_units = "Kelvin";

    pism_config:energy.temperature_based = "no";
    pism_config:energy.temperature_based_doc = "Use cold ice (i.e. not polythermal) methods.";
    pism_config:energy.temperature_based_type = "flag";

    pism_config:energy.temperature_dependent_thermal_conductivity = "no";
    pism_config:energy.temperature_dependent_thermal_conductivity_doc = "If yes, use varkenthSystemCtx class in the energy step. It is base on formula (4.37) in :cite:`GreveBlatter2009`. Otherwise use enthSystemCtx, which has temperature-independent thermal conductivity set by constant ice.thermal_conductivity.";
    pism_config:energy.temperature_dependent_thermal_conductivity_option = "vark";
    pism_config:energy.temperature_dependent_thermal_conductivity_type = "flag";

    pism_config:enthalpy_converter.T_reference = 223.15;
    pism_config:enthalpy_converter.T_reference_doc = "= T_0 in enthalpy formulas in :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_config:enthalpy_converter.T_reference_type = "number";
    pism_config:enthalpy_converter.T_reference_units = "Kelvin";

    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance = 0.001;
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_doc = "Tolerance within which ice is treated as temperate (cold-ice mode and diagnostics).";
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_type = "number";
    pism_config:enthalpy_converter.relaxed_is_temperate_tolerance_units = "Kelvin";

    pism_config:flow_law.Hooke.A = 4.42165e-9;
    pism_config:flow_law.Hooke.A_doc = "`A_{\\text{Hooke}} = (1/B_0)^n` where n=3 and `B_0` = 1.928 `a^{1/3}` Pa. See :cite:`Hooke`";
    pism_config:flow_law.Hooke.A_type = "number";
    pism_config:flow_law.Hooke.A_units = "Pascal-3 second-1";

    pism_config:flow_law.Hooke.C = 0.16612;
    pism_config:flow_law.Hooke.C_doc = "See :cite:`Hooke`";
    pism_config:flow_law.Hooke.C_type = "number";
    pism_config:flow_law.Hooke.C_units = "Kelvin^k";

    pism_config:flow_law.Hooke.Q = 7.88e4;
    pism_config:flow_law.Hooke.Q_doc = "Activation energy, see :cite:`Hooke`";
    pism_config:flow_law.Hooke.Q_type = "number";
    pism_config:flow_law.Hooke.Q_units = "Joule / mol";

    pism_config:flow_law.Hooke.Tr = 273.39;
    pism_config:flow_law.Hooke.Tr_doc = "See :cite:`Hooke`";
    pism_config:flow_law.Hooke.Tr_type = "number";
    pism_config:flow_law.Hooke.Tr_units = "Kelvin";

    pism_config:flow_law.Hooke.k = 1.17;
    pism_config:flow_law.Hooke.k_doc = "See :cite:`Hooke`";
    pism_config:flow_law.Hooke.k_type = "number";
    pism_config:flow_law.Hooke.k_units = "pure number";

    pism_config:flow_law.Paterson_Budd.A_cold = 3.61e-13;
    pism_config:flow_law.Paterson_Budd.A_cold_doc = "Paterson-Budd `A_\\text{cold}`, see :cite:`PatersonBudd`";
    pism_config:flow_law.Paterson_Budd.A_cold_type = "number";
    pism_config:flow_law.Paterson_Budd.A_cold_units = "Pascal-3 / second";

    pism_config:flow_law.Paterson_Budd.A_warm = 1.73e3;
    pism_config:flow_law.Paterson_Budd.A_warm_doc = "Paterson-Budd `A_\\text{warm}`, see :cite:`PatersonBudd`";
    pism_config:flow_law.Paterson_Budd.A_warm_type = "number";
    pism_config:flow_law.Paterson_Budd.A_warm_units = "Pascal-3 / second";

    pism_config:flow_law.Paterson_Budd.Q_cold = 6.0e4;
    pism_config:flow_law.Paterson_Budd.Q_cold_doc = "Paterson-Budd `Q_\\text{cold}`, see :cite:`PatersonBudd`";
    pism_config:flow_law.Paterson_Budd.Q_cold_type = "number";
    pism_config:flow_law.Paterson_Budd.Q_cold_units = "Joule / mol";

    pism_config:flow_law.Paterson_Budd.Q_warm = 13.9e4;
    pism_config:flow_law.Paterson_Budd.Q_warm_doc = "Paterson-Budd `Q_\\text{warm}`, see :cite:`PatersonBudd`";
    pism_config:flow_law.Paterson_Budd.Q_warm_type = "number";
    pism_config:flow_law.Paterson_Budd.Q_warm_units = "Joule / mol";

    pism_config:flow_law.Paterson_Budd.T_critical = 263.15;
    pism_config:flow_law.Paterson_Budd.T_critical_doc = "Paterson-Budd critical temperature, see :cite:`PatersonBudd`";
    pism_config:flow_law.Paterson_Budd.T_critical_type = "number";
    pism_config:flow_law.Paterson_Budd.T_critical_units = "Kelvin";

    pism_config:flow_law.Schoof_regularizing_length = 1000.0;
    pism_config:flow_law.Schoof_regularizing_length_doc = "Regularizing length (Schoof definition)";
    pism_config:flow_law.Schoof_regularizing_length_type = "number";
    pism_config:flow_law.Schoof_regularizing_length_units = "km";

    pism_config:flow_law.Schoof_regularizing_velocity = 1.0;
    pism_config:flow_law.Schoof_regularizing_velocity_doc = "Regularizing velocity (Schoof definition)";
    pism_config:flow_law.Schoof_regularizing_velocity_type = "number";
    pism_config:flow_law.Schoof_regularizing_velocity_units = "meter / year";

    pism_config:flow_law.gpbld.water_frac_coeff = 181.25;
    pism_config:flow_law.gpbld.water_frac_coeff_doc = "coefficient in Glen-Paterson-Budd flow law for extra dependence of softness on liquid water fraction (omega) :cite:`GreveBlatter2009`, :cite:`LliboutryDuval1985`";
    pism_config:flow_law.gpbld.water_frac_coeff_type = "number";
    pism_config:flow_law.gpbld.water_frac_coeff_units = "pure number";

    pism_config:flow_law.gpbld.water_frac_observed_limit = 0.01;
    pism_config:flow_law.gpbld.water_frac_observed_limit_doc = "maximum value of liquid water fraction omega for which softness values are parameterized by :cite:`LliboutryDuval1985`; used in Glen-Paterson-Budd-Lliboutry-Duval flow law; compare :cite:`AschwandenBuelerKhroulevBlatter`";
    pism_config:flow_law.gpbld.water_frac_observed_limit_type = "number";
    pism_config:flow_law.gpbld.water_frac_observed_limit_units = "1";

    pism_config:flow_law.isothermal_Glen.ice_softness = 3.1689e-24;
    pism_config:flow_law.isothermal_Glen.ice_softness_doc = "ice softness used by the isothermal Glen flow law :cite:`EISMINT96`";
    pism_config:flow_law.isothermal_Glen.ice_softness_type = "number";
    pism_config:flow_law.isothermal_Glen.ice_softness_units = "Pascal-3 second-1";

    pism_config:fracture_density.borstad_limit = "no";
    pism_config:fracture_density.borstad_limit_doc = "Model fracture growth according to the constitutive law in :cite:`Borstad2016Constitutive` (Eq. 4), ignoring :config:`fracture_density.gamma`.";
    pism_config:fracture_density.borstad_limit_option = "constitutive_stress_limit";
    pism_config:fracture_density.borstad_limit_type = "flag";

    pism_config:fracture_density.constant_fd = "no";
    pism_config:fracture_density.constant_fd_doc = "Keep fracture density fields constant in time but include its softening effect.";
    pism_config:fracture_density.constant_fd_option = "constant_fd";
    pism_config:fracture_density.constant_fd_type = "flag";

    pism_config:fracture_density.constant_healing = "no";
    pism_config:fracture_density.constant_healing_doc = "Use a constant healing rate `-\\gamma_h \\dot{\\epsilon}_h` independent of the local strain rate.";
    pism_config:fracture_density.constant_healing_option = "constant_healing";
    pism_config:fracture_density.constant_healing_type = "flag";

    pism_config:fracture_density.enabled = "no";
    pism_config:fracture_density.enabled_doc = "Model the fracture density using computed to stresses and strain rates.";
    pism_config:fracture_density.enabled_option = "fractures";
    pism_config:fracture_density.enabled_type = "flag";

    pism_config:fracture_density.fd2d_scheme = "no";
    pism_config:fracture_density.fd2d_scheme_doc = "Use an alternative transport scheme to reduce numerical diffusion (Eq. 10 in :cite:`AlbrechtLevermann2014softening`)";
    pism_config:fracture_density.fd2d_scheme_option = "scheme_fd2d";
    pism_config:fracture_density.fd2d_scheme_type = "flag";

    pism_config:fracture_density.fracture_weighted_healing = "no";
    pism_config:fracture_density.fracture_weighted_healing_doc = "Multiply the healing rate by `1 - D`, i.e. assume that highly damaged ice heals slower. This mechanism can be combined with :config:`fracture_density.constant_healing`.";
    pism_config:fracture_density.fracture_weighted_healing_option = "fracture_weighted_healing";
    pism_config:fracture_density.fracture_weighted_healing_type = "flag";

    pism_config:fracture_density.gamma = 1.0;
    pism_config:fracture_density.gamma_doc = "fracture growth constant `\\gamma`";
    pism_config:fracture_density.gamma_option = "fracture_gamma";
    pism_config:fracture_density.gamma_units = "1";
    pism_config:fracture_density.gamma_type = "number";

    pism_config:fracture_density.gamma_h = 0.0;
    pism_config:fracture_density.gamma_h_doc = "fracture healing constant `\\gamma_{h}`";
    pism_config:fracture_density.gamma_h_option = "fracture_gamma_h";
    pism_config:fracture_density.gamma_h_units = "1";
    pism_config:fracture_density.gamma_h_type = "number";

    pism_config:fracture_density.healing_threshold = 2.0e-10;
    pism_config:fracture_density.healing_threshold_doc = "fracture healing strain rate threshold `\\dot \\epsilon_{h}`";
    pism_config:fracture_density.healing_threshold_option = "fracture_healing_threshold";
    pism_config:fracture_density.healing_threshold_units = "1/s";
    pism_config:fracture_density.healing_threshold_type = "number";

    pism_config:fracture_density.include_grounded_ice = "no";
    pism_config:fracture_density.include_grounded_ice_doc = "Model fracture density in grounded areas (e.g. along ice stream shear zones) in addition to ice shelves";
    pism_config:fracture_density.include_grounded_ice_option = "do_frac_on_grounded";
    pism_config:fracture_density.include_grounded_ice_type = "flag";

    pism_config:fracture_density.initiation_threshold = 7.0e4;
    pism_config:fracture_density.initiation_threshold_doc = "fracture initiation stress threshold `\\sigma_{\\text{cr}}`";
    pism_config:fracture_density.initiation_threshold_option = "fracture_initiation_threshold";
    pism_config:fracture_density.initiation_threshold_units = "Pa";
    pism_config:fracture_density.initiation_threshold_type = "number";

    pism_config:fracture_density.lefm = "no";
    pism_config:fracture_density.lefm_doc = "Use the mixed-mode fracture toughness stress criterion based on Linear Elastic Fracture Mechanics, Eqs. 8-9 in :cite:`AlbrechtLevermann2014softening`";
    pism_config:fracture_density.lefm_option = "lefm";
    pism_config:fracture_density.lefm_type = "flag";

    pism_config:fracture_density.max_shear_stress = "no";
    pism_config:fracture_density.max_shear_stress_doc = "Use the maximum shear stress criterion for fracture formation (Tresca or Guest criterion in literature), which is more stringent than the default von Mises criterion, see Eq. 7 in :cite:`AlbrechtLevermann2014softening`";
    pism_config:fracture_density.max_shear_stress_option = "max_shear";
    pism_config:fracture_density.max_shear_stress_type = "flag";

    pism_config:fracture_density.phi0 = 0.0;
    pism_config:fracture_density.phi0_doc = "Fracture density value used at grid points where ice velocity is prescribed. This assumes that all ice entering a shelf at :var:`bc_mask` locations has the same fracture density.";
    pism_config:fracture_density.phi0_option = "phi0";
    pism_config:fracture_density.phi0_type = "number";
    pism_config:fracture_density.phi0_units = "1";

    pism_config:fracture_density.softening_lower_limit = 1.0;
    pism_config:fracture_density.softening_lower_limit_doc = "Parameter controlling the strength of the feedback of damage on the ice flow. If `1`: no feedback, if `0`: full feedback (`\\epsilon` in Eq. 6 in :cite:`AlbrechtLevermann2014softening`)";
    pism_config:fracture_density.softening_lower_limit_option = "fracture_softening";
    pism_config:fracture_density.softening_lower_limit_type = "number";
    pism_config:fracture_density.softening_lower_limit_units = "1";

    pism_config:frontal_melt.constant.melt_rate = 1.0;
    pism_config:frontal_melt.constant.melt_rate_doc = "default melt rate used by the ``constant`` frontal_melt model";
    pism_config:frontal_melt.constant.melt_rate_option = "frontal_melt_rate";
    pism_config:frontal_melt.constant.melt_rate_type = "number";
    pism_config:frontal_melt.constant.melt_rate_units = "m / day";

    pism_config:frontal_melt.discharge_given.file = "";
    pism_config:frontal_melt.discharge_given.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:frontal_melt.discharge_given.file_option = "frontal_melt_discharge_given_file";
    pism_config:frontal_melt.discharge_given.file_type = "string";

    pism_config:frontal_melt.discharge_given.periodic = "no";
    pism_config:frontal_melt.discharge_given.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:frontal_melt.discharge_given.periodic_type = "flag";

    pism_config:frontal_melt.given.file = "";
    pism_config:frontal_melt.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:frontal_melt.given.file_option = "frontal_melt_given_file";
    pism_config:frontal_melt.given.file_type = "string";

    pism_config:frontal_melt.given.periodic = "no";
    pism_config:frontal_melt.given.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:frontal_melt.given.periodic_type = "flag";

    pism_config:frontal_melt.include_floating_ice = "no";
    pism_config:frontal_melt.include_floating_ice_doc = "Apply frontal melt to all grid icy cells next to ocean cells";
    pism_config:frontal_melt.include_floating_ice_type = "flag";

    pism_config:frontal_melt.models = "";
    pism_config:frontal_melt.models_doc = "Comma-separated list of frontal melt models and modifiers. (Leave empty to disable.)";
    pism_config:frontal_melt.models_option = "frontal_melt";
    pism_config:frontal_melt.models_type = "string";

    pism_config:frontal_melt.open_ocean_margins_only = "no";
    pism_config:frontal_melt.open_ocean_margins_only_doc = "Apply frontal melt parameterizations only at ice fronts bordering ice-free ocean areas that are connected to the open ocean";
    pism_config:frontal_melt.open_ocean_margins_only_type = "flag";

    pism_config:frontal_melt.routing.file = "";
    pism_config:frontal_melt.routing.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:frontal_melt.routing.file_option = "frontal_melt_routing_file";
    pism_config:frontal_melt.routing.file_type = "string";

    pism_config:frontal_melt.routing.parameter_a = 3e-4;
    pism_config:frontal_melt.routing.parameter_a_doc = "parameter A in eqn. 1 in :cite:`Xu2013`";
    pism_config:frontal_melt.routing.parameter_a_type = "number";
    pism_config:frontal_melt.routing.parameter_a_units = "m-alpha day^(alpha-1) Celsius-beta";

    pism_config:frontal_melt.routing.parameter_b = 0.15;
    pism_config:frontal_melt.routing.parameter_b_doc = "parameter B in eqn. 1 in :cite:`Xu2013`";
    pism_config:frontal_melt.routing.parameter_b_type = "number";
    pism_config:frontal_melt.routing.parameter_b_units = "m day^(alpha-1) Celsius-beta";

    pism_config:frontal_melt.routing.periodic = "no";
    pism_config:frontal_melt.routing.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:frontal_melt.routing.periodic_type = "flag";

    pism_config:frontal_melt.routing.power_alpha = 0.39;
    pism_config:frontal_melt.routing.power_alpha_doc = "exponent `\\alpha` in eqn. 1 in :cite:`Xu2013`";
    pism_config:frontal_melt.routing.power_alpha_type = "number";
    pism_config:frontal_melt.routing.power_alpha_units = "1";

    pism_config:frontal_melt.routing.power_beta = 1.18;
    pism_config:frontal_melt.routing.power_beta_doc = "exponent `\\beta` in eqn. 1 in :cite:`Xu2013`";
    pism_config:frontal_melt.routing.power_beta_type = "number";
    pism_config:frontal_melt.routing.power_beta_units = "1";

    pism_config:geometry.front_retreat.minimum_time_step = 0.01;
    pism_config:geometry.front_retreat.minimum_time_step_doc = "Minimum allowed time step length. Increase this to keep calving models from slowing PISM down too much.";
    pism_config:geometry.front_retreat.minimum_time_step_units = "365day";
    pism_config:geometry.front_retreat.minimum_time_step_type = "number";

    pism_config:geometry.front_retreat.prescribed.file = "";
    pism_config:geometry.front_retreat.prescribed.file_doc = "Name of the file containing the maximum ice extent mask ``land_ice_area_fraction_retreat``";
    pism_config:geometry.front_retreat.prescribed.file_option = "front_retreat_file";
    pism_config:geometry.front_retreat.prescribed.file_type = "string";

    pism_config:geometry.front_retreat.prescribed.periodic = "no";
    pism_config:geometry.front_retreat.prescribed.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:geometry.front_retreat.prescribed.periodic_type = "flag";

    pism_config:geometry.front_retreat.use_cfl = "false";
    pism_config:geometry.front_retreat.use_cfl_doc = "apply CFL criterion for eigen-calving rate front retreat";
    pism_config:geometry.front_retreat.use_cfl_option = "front_retreat_cfl";
    pism_config:geometry.front_retreat.use_cfl_type = "flag";

    pism_config:geometry.front_retreat.wrap_around = "false";
    pism_config:geometry.front_retreat.wrap_around_doc = "If true, wrap around domain boundaries. This may be needed in some regional synthetic geometry setups.";
    pism_config:geometry.front_retreat.wrap_around_option = "front_retreat_wrap_around";
    pism_config:geometry.front_retreat.wrap_around_type = "flag";

    pism_config:geometry.grounded_cell_fraction  = "false";
    pism_config:geometry.grounded_cell_fraction_doc = "Linear interpolation scheme (\"LI\" in Gladstone et al. 2010) expanded to two dimensions is used if switched on in order to evaluate the position of the grounding line on a subgrid scale.";
    pism_config:geometry.grounded_cell_fraction_option = "subgl";
    pism_config:geometry.grounded_cell_fraction_type = "flag";

    pism_config:geometry.ice_free_thickness_standard = 0.01;
    pism_config:geometry.ice_free_thickness_standard_doc = "If ice is thinner than this standard then the mask is set to MASK_ICE_FREE_BEDROCK or MASK_ICE_FREE_OCEAN.";
    pism_config:geometry.ice_free_thickness_standard_type = "number";
    pism_config:geometry.ice_free_thickness_standard_units = "meters";

    pism_config:geometry.part_grid.enabled = "no";
    pism_config:geometry.part_grid.enabled_doc = "apply partially filled grid cell scheme";
    pism_config:geometry.part_grid.enabled_option = "part_grid";
    pism_config:geometry.part_grid.enabled_type = "flag";

    pism_config:geometry.part_grid.max_iterations = 10;
    pism_config:geometry.part_grid.max_iterations_doc = "maximum number of residual redistribution iterations";
    pism_config:geometry.part_grid.max_iterations_type = "integer";
    pism_config:geometry.part_grid.max_iterations_units = "count";

    pism_config:geometry.remove_icebergs = "no";
    pism_config:geometry.remove_icebergs_doc = "identify and kill detached ice-shelf areas";
    pism_config:geometry.remove_icebergs_option = "kill_icebergs";
    pism_config:geometry.remove_icebergs_type = "flag";

    pism_config:geometry.update.enabled = "yes";
    pism_config:geometry.update.enabled_doc = "Solve the mass conservation equation";
    pism_config:geometry.update.enabled_option = "mass";
    pism_config:geometry.update.enabled_type = "flag";

    pism_config:geometry.update.use_basal_melt_rate = "yes";
    pism_config:geometry.update.use_basal_melt_rate_doc = "Include basal melt rate in the continuity equation";
    pism_config:geometry.update.use_basal_melt_rate_option = "bmr_in_cont";
    pism_config:geometry.update.use_basal_melt_rate_type = "flag";

    pism_config:grid.Lbz = 1000;
    pism_config:grid.Lbz_doc = "Thickness of the thermal bedrock layer. (Inactive if :config:`grid.Mbz` < 2)";
    pism_config:grid.Lbz_option = "Lbz";
    pism_config:grid.Lbz_type = "number";
    pism_config:grid.Lbz_units = "meters";

    pism_config:grid.Lx = 1500e3;
    pism_config:grid.Lx_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_config:grid.Lx_type = "number";
    pism_config:grid.Lx_units = "meters";

    pism_config:grid.Ly = 1500e3;
    pism_config:grid.Ly_doc = "Default computational box is 3000 km x 3000 km (= 2 Lx x 2 Ly) in horizontal.";
    pism_config:grid.Ly_type = "number";
    pism_config:grid.Ly_units = "meters";

    pism_config:grid.Lz = 4000;
    pism_config:grid.Lz_doc = "Height of the computational domain.";
    pism_config:grid.Lz_option = "Lz";
    pism_config:grid.Lz_type = "number";
    pism_config:grid.Lz_units = "meters";

    pism_config:grid.Mbz = 1;
    pism_config:grid.Mbz_doc = "Number of thermal bedrock layers; 1 level corresponds to no bedrock.";
    pism_config:grid.Mbz_option = "Mbz";
    pism_config:grid.Mbz_type = "integer";
    pism_config:grid.Mbz_units = "count";

    pism_config:grid.Mx = 61;
    pism_config:grid.Mx_doc = "Number of grid points in the x direction.";
    pism_config:grid.Mx_option = "Mx";
    pism_config:grid.Mx_type = "integer";
    pism_config:grid.Mx_units = "count";

    pism_config:grid.My = 61;
    pism_config:grid.My_doc = "Number of grid points in the y direction.";
    pism_config:grid.My_option = "My";
    pism_config:grid.My_type = "integer";
    pism_config:grid.My_units = "count";

    pism_config:grid.Mz = 31;
    pism_config:grid.Mz_doc = "Number of vertical grid levels in the ice.";
    pism_config:grid.Mz_option = "Mz";
    pism_config:grid.Mz_type = "integer";
    pism_config:grid.Mz_units = "count";

    pism_config:grid.allow_extrapolation = "no";
    pism_config:grid.allow_extrapolation_doc = "Allow extrapolation during regridding.";
    pism_config:grid.allow_extrapolation_option = "allow_extrapolation";
    pism_config:grid.allow_extrapolation_type = "flag";

    pism_config:grid.ice_vertical_spacing = "quadratic";
    pism_config:grid.ice_vertical_spacing_choices = "quadratic,equal";
    pism_config:grid.ice_vertical_spacing_doc = "vertical spacing in the ice";
    pism_config:grid.ice_vertical_spacing_option = "z_spacing";
    pism_config:grid.ice_vertical_spacing_type = "keyword";

    pism_config:grid.lambda = 4.0;
    pism_config:grid.lambda_doc = "Vertical grid spacing parameter. Roughly equal to the factor by which the grid is coarser at an end away from the ice-bedrock interface.";
    pism_config:grid.lambda_type = "number";
    pism_config:grid.lambda_units = "pure number";

    pism_config:grid.max_stencil_width = 2;
    pism_config:grid.max_stencil_width_doc = "Maximum width of the finite-difference stencil used in PISM.";
    pism_config:grid.max_stencil_width_type = "integer";
    pism_config:grid.max_stencil_width_units = "count";

    pism_config:grid.periodicity = "xy";
    pism_config:grid.periodicity_choices = "none,x,y,xy";
    pism_config:grid.periodicity_doc = "horizontal grid periodicity";
    pism_config:grid.periodicity_option = "periodicity";
    pism_config:grid.periodicity_type = "keyword";

    pism_config:grid.recompute_longitude_and_latitude = "yes";
    pism_config:grid.recompute_longitude_and_latitude_doc = "Re-compute longitude and latitude using grid information and provided projection parameters. Requires PROJ.";
    pism_config:grid.recompute_longitude_and_latitude_type = "flag";

    pism_config:grid.registration = "center";
    pism_config:grid.registration_choices = "center,corner";
    pism_config:grid.registration_doc = "horizontal grid registration";
    pism_config:grid.registration_type = "keyword";

    pism_config:hydrology.add_water_input_to_till_storage = "yes";
    pism_config:hydrology.add_water_input_to_till_storage_doc = "Add surface input to water stored in till. If no it will be added to the transportable water.";
    pism_config:hydrology.add_water_input_to_till_storage_type = "flag";

    pism_config:hydrology.cavitation_opening_coefficient = 0.5;
    pism_config:hydrology.cavitation_opening_coefficient_doc = "c_1 in notes; coefficient of cavitation opening term in evolution of layer thickness in hydrology::Distributed";
    pism_config:hydrology.cavitation_opening_coefficient_option = "hydrology_cavitation_opening_coefficient";
    pism_config:hydrology.cavitation_opening_coefficient_type = "number";
    pism_config:hydrology.cavitation_opening_coefficient_units = "meter-1";

    pism_config:hydrology.creep_closure_coefficient = 0.04;
    pism_config:hydrology.creep_closure_coefficient_doc = "c_2 in notes; coefficient of creep closure term in evolution of layer thickness in hydrology::Distributed";
    pism_config:hydrology.creep_closure_coefficient_option = "hydrology_creep_closure_coefficient";
    pism_config:hydrology.creep_closure_coefficient_type = "number";
    pism_config:hydrology.creep_closure_coefficient_units = "pure number";

    pism_config:hydrology.distributed.init_p_from_steady = "no";
    pism_config:hydrology.distributed.init_p_from_steady_doc = "if \"yes\", initialize subglacial water pressure from P(W) formula that applies in steady state";
    pism_config:hydrology.distributed.init_p_from_steady_option = "hydrology_init_p_form_steady";
    pism_config:hydrology.distributed.init_p_from_steady_type = "flag";

    pism_config:hydrology.distributed.sliding_speed_file = "";
    pism_config:hydrology.distributed.sliding_speed_file_doc = "name of the file containing velbase_mag, the basal sliding speed to use with :literal:`hydrology.distributed.init_p_from_steady`";
    pism_config:hydrology.distributed.sliding_speed_file_option = "hydrology_sliding_speed_file";
    pism_config:hydrology.distributed.sliding_speed_file_type = "string";

    pism_config:hydrology.gradient_power_in_flux = 1.5;
    pism_config:hydrology.gradient_power_in_flux_doc = "power `\\beta` in Darcy's law `q = - k W^{\\alpha} |\\nabla \\psi|^{\\beta-2} \\nabla \\psi`, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.gradient_power_in_flux_option = "hydrology_gradient_power_in_flux";
    pism_config:hydrology.gradient_power_in_flux_type = "number";
    pism_config:hydrology.gradient_power_in_flux_units = "pure number";

    pism_config:hydrology.hydraulic_conductivity = 0.001;
    pism_config:hydrology.hydraulic_conductivity_doc = "= k in notes; lateral conductivity, in Darcy's law, for subglacial water layer; units depend on powers alpha = hydrology.thickness_power_in_flux and beta = hydrology_potential_gradient_power_in_flux; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.hydraulic_conductivity_option = "hydrology_hydraulic_conductivity";
    pism_config:hydrology.hydraulic_conductivity_type = "number";
    pism_config:hydrology.hydraulic_conductivity_units = "`m^{2 \\beta - \\alpha} s^{2 \\beta - 3} kg^{1-\\beta}`";

    pism_config:hydrology.maximum_time_step = 1.0;
    pism_config:hydrology.maximum_time_step_doc = "maximum allowed time step length used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.maximum_time_step_type = "number";
    pism_config:hydrology.maximum_time_step_units = "365days";

    pism_config:hydrology.model = "null";
    pism_config:hydrology.model_choices = "null,routing,steady,distributed";
    pism_config:hydrology.model_doc = "Basal hydrology sub-model.";
    pism_config:hydrology.model_option = "hydrology";
    pism_config:hydrology.model_type = "keyword";

    pism_config:hydrology.null_diffuse_till_water = "no";
    pism_config:hydrology.null_diffuse_till_water_doc = "Diffuse stored till water laterally. See equation (11) of :cite:`BBssasliding`";
    pism_config:hydrology.null_diffuse_till_water_type = "flag";

    pism_config:hydrology.null_diffusion_distance = 2e4;
    pism_config:hydrology.null_diffusion_distance_doc = "diffusion distance for till water thickness; see equation (11) in :cite:`BBssasliding`; only active if hydrology.null_diffuse_till_water is set";
    pism_config:hydrology.null_diffusion_distance_type = "number";
    pism_config:hydrology.null_diffusion_distance_units = "meters";

    pism_config:hydrology.null_diffusion_time = 1000.0;
    pism_config:hydrology.null_diffusion_time_doc = "diffusion time for till water thickness; see equation (11) in :cite:`BBssasliding`; only active if hydrology.null_diffuse_till_water is set";
    pism_config:hydrology.null_diffusion_time_type = "number";
    pism_config:hydrology.null_diffusion_time_units = "365days";

    pism_config:hydrology.regularizing_porosity = 0.01;
    pism_config:hydrology.regularizing_porosity_doc = "phi_0 in notes; regularizes pressure equation by multiplying time derivative term";
    pism_config:hydrology.regularizing_porosity_option = "hydrology_regularizing_porosity";
    pism_config:hydrology.regularizing_porosity_type = "number";
    pism_config:hydrology.regularizing_porosity_units = "pure number";

    pism_config:hydrology.roughness_scale = 0.1;
    pism_config:hydrology.roughness_scale_doc = "W_r in notes; roughness scale determining maximum amount of cavitation opening in hydrology::Distributed";
    pism_config:hydrology.roughness_scale_option = "hydrology_roughness_scale";
    pism_config:hydrology.roughness_scale_type = "number";
    pism_config:hydrology.roughness_scale_units = "meters";

    pism_config:hydrology.routing.include_floating_ice = "no";
    pism_config:hydrology.routing.include_floating_ice_doc = "Route subglacial water under ice shelves. This may be appropriate if a shelf is close to floatation. Note that this has no effect on ice flow.";
    pism_config:hydrology.routing.include_floating_ice_type = "flag";

    pism_config:hydrology.steady.flux_update_interval = 1.0;
    pism_config:hydrology.steady.flux_update_interval_doc = "interval between updates of the steady state flux";
    pism_config:hydrology.steady.flux_update_interval_type = "number";
    pism_config:hydrology.steady.flux_update_interval_units = "365days";

    pism_config:hydrology.steady.input_rate_scaling = 1e7;
    pism_config:hydrology.steady.input_rate_scaling_doc = "input rate scaling";
    pism_config:hydrology.steady.input_rate_scaling_type = "number";
    pism_config:hydrology.steady.input_rate_scaling_units = "seconds";

    pism_config:hydrology.steady.n_iterations = 7500;
    pism_config:hydrology.steady.n_iterations_doc = "maxinum number of iterations to use in while estimating steady-state water flux";
    pism_config:hydrology.steady.n_iterations_type = "integer";
    pism_config:hydrology.steady.n_iterations_units = "count";

    pism_config:hydrology.steady.potential_delta = 10000.0;
    pism_config:hydrology.steady.potential_delta_doc = "potential adjustment used to fill sinks (smaller values require more iterations but produce fewer artifacts)";
    pism_config:hydrology.steady.potential_delta_type = "number";
    pism_config:hydrology.steady.potential_delta_units = "Pa";

    pism_config:hydrology.steady.potential_n_iterations = 1000;
    pism_config:hydrology.steady.potential_n_iterations_doc = "maxinum number of iterations to take while pre-processing hydraulic potential";
    pism_config:hydrology.steady.potential_n_iterations_type = "integer";
    pism_config:hydrology.steady.potential_n_iterations_units = "count";

    pism_config:hydrology.steady.volume_ratio = 0.1;
    pism_config:hydrology.steady.volume_ratio_doc = "water volume ratio used as the stopping criterion";
    pism_config:hydrology.steady.volume_ratio_type = "number";
    pism_config:hydrology.steady.volume_ratio_units = "1";

    pism_config:hydrology.surface_input.file = "";
    pism_config:hydrology.surface_input.file_doc = "Name of the file containing :var:`water_input_rate`, the rate at which water from the ice surface is added to the subglacial hydrology system";
    pism_config:hydrology.surface_input.file_type = "string";

    pism_config:hydrology.surface_input.periodic = "no";
    pism_config:hydrology.surface_input.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:hydrology.surface_input.periodic_type = "flag";

    pism_config:hydrology.surface_input_from_runoff = "no";
    pism_config:hydrology.surface_input_from_runoff_doc = "Use surface runoff as surface input.";
    pism_config:hydrology.surface_input_from_runoff_type = "flag";

    pism_config:hydrology.thickness_power_in_flux = 1.25;
    pism_config:hydrology.thickness_power_in_flux_doc = "power `\\alpha` in Darcy's law `q = - k W^{\\alpha} |\\nabla \\psi|^{\\beta-2} \\nabla \\psi`, for subglacial water layer; used by hydrology::Routing and hydrology::Distributed";
    pism_config:hydrology.thickness_power_in_flux_option = "hydrology_thickness_power_in_flux";
    pism_config:hydrology.thickness_power_in_flux_type = "number";
    pism_config:hydrology.thickness_power_in_flux_units = "1";

    pism_config:hydrology.tillwat_decay_rate = 1.0;
    pism_config:hydrology.tillwat_decay_rate_doc = "rate at which tillwat is reduced to zero, in absence of other effects like input";
    pism_config:hydrology.tillwat_decay_rate_option = "hydrology_tillwat_decay_rate";
    pism_config:hydrology.tillwat_decay_rate_type = "number";
    pism_config:hydrology.tillwat_decay_rate_units = "mm / year";

    pism_config:hydrology.tillwat_max = 2.0;
    pism_config:hydrology.tillwat_max_doc = "maximum effective thickness of the water stored in till";
    pism_config:hydrology.tillwat_max_option = "hydrology_tillwat_max";
    pism_config:hydrology.tillwat_max_type = "number";
    pism_config:hydrology.tillwat_max_units = "meters";

    pism_config:input.bootstrap = "no";
    pism_config:input.bootstrap_doc = "It true, use bootstrapping heuristics when initializing PISM.";
    pism_config:input.bootstrap_option = "bootstrap";
    pism_config:input.bootstrap_type = "flag";

    pism_config:input.file = "";
    pism_config:input.file_doc = "Input file name";
    pism_config:input.file_option = "i";
    pism_config:input.file_type = "string";

    pism_config:input.forcing.buffer_size = 60;
    pism_config:input.forcing.buffer_size_doc = "number of 2D climate forcing records to keep in memory; = 5 years of monthly records";
    pism_config:input.forcing.buffer_size_type = "integer";
    pism_config:input.forcing.buffer_size_units = "count";

    pism_config:input.forcing.time_extrapolation = "false";
    pism_config:input.forcing.time_extrapolation_doc = "If 'true', time-dependent forcing inputs are extrapolated in time";
    pism_config:input.forcing.time_extrapolation_type = "flag";

    pism_config:input.regrid.file = "";
    pism_config:input.regrid.file_doc = "Regridding (input) file name";
    pism_config:input.regrid.file_option = "regrid_file";
    pism_config:input.regrid.file_type = "string";

    pism_config:input.regrid.vars = "";
    pism_config:input.regrid.vars_doc = "Comma-separated list of variables to regrid. Leave empty to regrid all model state variables.";
    pism_config:input.regrid.vars_option = "regrid_vars";
    pism_config:input.regrid.vars_type = "string";

    pism_config:inverse.design.cH1     = 0;
    pism_config:inverse.design.cH1_doc = "weight of derivative part of an H1 norm for inversion design variables";
    pism_config:inverse.design.cH1_option = "inv_design_cH1";
    pism_config:inverse.design.cH1_type = "number";
    pism_config:inverse.design.cH1_units = "1";

    pism_config:inverse.design.cL2 = 1;
    pism_config:inverse.design.cL2_doc = "weight of derivative-free part of an H1 norm for inversion design variables";
    pism_config:inverse.design.cL2_option = "inv_design_cL2";
    pism_config:inverse.design.cL2_type = "number";
    pism_config:inverse.design.cL2_units = "1";

    pism_config:inverse.design.func = "sobolevH1";
    pism_config:inverse.design.func_choices = "sobolevH1,tv";
    pism_config:inverse.design.func_doc = "functional used for inversion design variables";
    pism_config:inverse.design.func_option = "inv_design_func";
    pism_config:inverse.design.func_type = "keyword";

    pism_config:inverse.design.param = "exp";
    pism_config:inverse.design.param_choices = "ident,trunc,square,exp";
    pism_config:inverse.design.param_doc = "parameterization of design variables used during inversion";
    pism_config:inverse.design.param_option = "inv_design_param";
    pism_config:inverse.design.param_type = "keyword";

    pism_config:inverse.design.param_tauc_eps = 100;
    pism_config:inverse.design.param_tauc_eps_doc = "tiny yield stress used as a substitute for 0 in some tauc parameterizations";
    pism_config:inverse.design.param_tauc_eps_type = "number";
    pism_config:inverse.design.param_tauc_eps_units = "Pascal";

    pism_config:inverse.design.param_tauc_scale = 100000;
    pism_config:inverse.design.param_tauc_scale_doc = "typical size of yield stresses";
    pism_config:inverse.design.param_tauc_scale_type = "number";
    pism_config:inverse.design.param_tauc_scale_units = "Pascal";

    pism_config:inverse.design.param_trunc_tauc0 = 1000;
    pism_config:inverse.design.param_trunc_tauc0_doc = "transition point of change to linear behaviour for design variable parameterization type ``trunc``";
    pism_config:inverse.design.param_trunc_tauc0_type = "number";
    pism_config:inverse.design.param_trunc_tauc0_units = "Pascal";

    pism_config:inverse.log_ratio_scale = 10;
    pism_config:inverse.log_ratio_scale_doc = "Reference scale for log-ratio functionals";
    pism_config:inverse.log_ratio_scale_option = "inv_log_ratio_scale";
    pism_config:inverse.log_ratio_scale_type = "number";
    pism_config:inverse.log_ratio_scale_units = "pure number";

    pism_config:inverse.max_iterations = 1000;
    pism_config:inverse.max_iterations_doc = "maximum iteration count";
    pism_config:inverse.max_iterations_option = "inv_max_it";
    pism_config:inverse.max_iterations_type = "integer";
    pism_config:inverse.max_iterations_units = "count";

    pism_config:inverse.ssa.hardav_max = 1e10;
    pism_config:inverse.ssa.hardav_max_doc = "Maximum allowed value of hardav for inversions with bound constraints";
    pism_config:inverse.ssa.hardav_max_type = "number";
    pism_config:inverse.ssa.hardav_max_units = "Pascal second^(1/3)";

    pism_config:inverse.ssa.hardav_min = 0;
    pism_config:inverse.ssa.hardav_min_doc = "Minimum allowed value of hardav for inversions with bound constraints";
    pism_config:inverse.ssa.hardav_min_type = "number";
    pism_config:inverse.ssa.hardav_min_units = "Pascal second^(1/3)";

    pism_config:inverse.ssa.length_scale = 50e3;
    pism_config:inverse.ssa.length_scale_doc = "typical length scale for rescaling derivative norms";
    pism_config:inverse.ssa.length_scale_type = "number";
    pism_config:inverse.ssa.length_scale_units = "meters";

    pism_config:inverse.ssa.method = "tikhonov_lmvm";
    pism_config:inverse.ssa.method_choices = "sd,nlcg,ign,tikhonov_lmvm,tikhonov_cg,tikhonov_blmvm,tikhonov_lcl,tikhonov_gn";
    pism_config:inverse.ssa.method_doc = "algorithm to use for SSA inversions";
    pism_config:inverse.ssa.method_option = "inv_method";
    pism_config:inverse.ssa.method_type = "keyword";

    pism_config:inverse.ssa.tauc_max = 5e7;
    pism_config:inverse.ssa.tauc_max_doc = "Maximum allowed value of tauc for inversions with bound constraints";
    pism_config:inverse.ssa.tauc_max_type = "number";
    pism_config:inverse.ssa.tauc_max_units = "Pascal";

    pism_config:inverse.ssa.tauc_min = 0;
    pism_config:inverse.ssa.tauc_min_doc = "Minimum allowed value of tauc for inversions with bound constraints";
    pism_config:inverse.ssa.tauc_min_type = "number";
    pism_config:inverse.ssa.tauc_min_units = "Pascal";

    pism_config:inverse.ssa.tv_exponent = 1.2;
    pism_config:inverse.ssa.tv_exponent_doc = "Lebesgue exponent for pseudo-TV norm";
    pism_config:inverse.ssa.tv_exponent_option = "inv_ssa_tv_exponent";
    pism_config:inverse.ssa.tv_exponent_type = "number";
    pism_config:inverse.ssa.tv_exponent_units = "pure number";

    pism_config:inverse.ssa.velocity_eps = 0.1;
    pism_config:inverse.ssa.velocity_eps_doc = "tiny size of ice velocities during inversion";
    pism_config:inverse.ssa.velocity_eps_type = "number";
    pism_config:inverse.ssa.velocity_eps_units = "meter / year";

    pism_config:inverse.ssa.velocity_scale = 100;
    pism_config:inverse.ssa.velocity_scale_doc = "typical size of ice velocities expected during inversion";
    pism_config:inverse.ssa.velocity_scale_type = "number";
    pism_config:inverse.ssa.velocity_scale_units = "meter / year";

    pism_config:inverse.state_func = "meansquare";
    pism_config:inverse.state_func_choices = "meansquare,log_ratio,log_relative";
    pism_config:inverse.state_func_doc = "functional used for inversion design variables";
    pism_config:inverse.state_func_option = "inv_state_func";
    pism_config:inverse.state_func_type = "keyword";

    pism_config:inverse.tikhonov.atol = 1e-10;
    pism_config:inverse.tikhonov.atol_doc = "absolute threshold for Tikhonov stopping criterion";
    pism_config:inverse.tikhonov.atol_option = "tikhonov_atol";
    pism_config:inverse.tikhonov.atol_type = "number";
    pism_config:inverse.tikhonov.atol_units = "meter / year";

    pism_config:inverse.tikhonov.penalty_weight = 1;
    pism_config:inverse.tikhonov.penalty_weight_doc = "penalty parameter for Tikhonov inversion";
    pism_config:inverse.tikhonov.penalty_weight_option = "tikhonov_penalty";
    pism_config:inverse.tikhonov.penalty_weight_type = "number";
    pism_config:inverse.tikhonov.penalty_weight_units = "1";

    pism_config:inverse.tikhonov.ptol = 0.1;
    pism_config:inverse.tikhonov.ptol_doc = "threshold for reaching desired misfit for adaptive Tikhonov algorithms";
    pism_config:inverse.tikhonov.ptol_option = "tikhonov_ptol";
    pism_config:inverse.tikhonov.ptol_type = "number";
    pism_config:inverse.tikhonov.ptol_units = "pure number";

    pism_config:inverse.tikhonov.rtol = 5e-2;
    pism_config:inverse.tikhonov.rtol_doc = "relative threshold for Tikhonov stopping criterion";
    pism_config:inverse.tikhonov.rtol_option = "tikhonov_rtol";
    pism_config:inverse.tikhonov.rtol_type = "number";
    pism_config:inverse.tikhonov.rtol_units = "1";

    pism_config:inverse.use_design_prior = "yes";
    pism_config:inverse.use_design_prior_doc = "Use prior from inverse data file as initial guess.";
    pism_config:inverse.use_design_prior_option = "inv_use_design_prior";
    pism_config:inverse.use_design_prior_type = "flag";

    pism_config:inverse.use_zeta_fixed_mask = "yes";
    pism_config:inverse.use_zeta_fixed_mask_doc = "Enforce locations where the parameterized design variable should be fixed. (Automatically determined if not provided)";
    pism_config:inverse.use_zeta_fixed_mask_option = "inv_use_zeta_fixed_mask";
    pism_config:inverse.use_zeta_fixed_mask_type = "flag";

    pism_config:isochrones.bootstrapping.n_layers = 0;
    pism_config:isochrones.bootstrapping.n_layers_doc = "number of isochronal layers created during bootstrapping";
    pism_config:isochrones.bootstrapping.n_layers_type = "integer";
    pism_config:isochrones.bootstrapping.n_layers_units = "count";

    pism_config:isochrones.deposition_times = "";
    pism_config:isochrones.deposition_times_doc = "List or a range of deposition times used to create isochronal layers";
    pism_config:isochrones.deposition_times_type = "string";

    pism_config:isochrones.max_n_layers = 100;
    pism_config:isochrones.max_n_layers_doc = "maximum number of isochronal layers";
    pism_config:isochrones.max_n_layers_type = "integer";
    pism_config:isochrones.max_n_layers_units = "count";

    pism_config:ocean.anomaly.file = "";
    pism_config:ocean.anomaly.file_doc = "Name of the file containing shelf basal mass flux offset fields.";
    pism_config:ocean.anomaly.file_option = "ocean_anomaly_file";
    pism_config:ocean.anomaly.file_type = "string";

    pism_config:ocean.anomaly.periodic = "no";
    pism_config:ocean.anomaly.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.anomaly.periodic_type = "flag";

    pism_config:ocean.cache.update_interval = 10;
    pism_config:ocean.cache.update_interval_doc = "update interval of the ``cache`` ocean modifier";
    pism_config:ocean.cache.update_interval_option = "ocean_cache_update_interval";
    pism_config:ocean.cache.update_interval_type = "integer";
    pism_config:ocean.cache.update_interval_units = "365days";

    pism_config:ocean.constant.melt_rate = 0.05191419359084029;
    pism_config:ocean.constant.melt_rate_doc = "default melt rate used by the ``constant`` ocean model (computed as `Q / (L \\rho_i)`)";
    pism_config:ocean.constant.melt_rate_option = "shelf_base_melt_rate";
    pism_config:ocean.constant.melt_rate_type = "number";
    pism_config:ocean.constant.melt_rate_units = "m / year";

    pism_config:ocean.delta_MBP.file = "";
    pism_config:ocean.delta_MBP.file_doc = "Name of the file containing melange back-pressure offsets";
    pism_config:ocean.delta_MBP.file_type = "string";

    pism_config:ocean.delta_MBP.melange_thickness = 100.0;
    pism_config:ocean.delta_MBP.melange_thickness_doc = "Melange thickness (assumed to be constant in space and time)";
    pism_config:ocean.delta_MBP.melange_thickness_option = "melange_thickness";
    pism_config:ocean.delta_MBP.melange_thickness_type = "number";
    pism_config:ocean.delta_MBP.melange_thickness_units = "meters";

    pism_config:ocean.delta_MBP.periodic = "no";
    pism_config:ocean.delta_MBP.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.delta_MBP.periodic_type = "flag";

    pism_config:ocean.delta_T.file = "";
    pism_config:ocean.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_config:ocean.delta_T.file_option = "ocean_delta_T_file";
    pism_config:ocean.delta_T.file_type = "string";

    pism_config:ocean.delta_T.periodic = "no";
    pism_config:ocean.delta_T.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.delta_T.periodic_type = "flag";

    pism_config:ocean.delta_mass_flux.file = "";
    pism_config:ocean.delta_mass_flux.file_doc = "Name of the file containing sub-shelf mass flux offsets.";
    pism_config:ocean.delta_mass_flux.file_option = "ocean_delta_mass_flux_file";
    pism_config:ocean.delta_mass_flux.file_type = "string";

    pism_config:ocean.delta_mass_flux.periodic = "no";
    pism_config:ocean.delta_mass_flux.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.delta_mass_flux.periodic_type = "flag";

    pism_config:ocean.delta_sl.file = "";
    pism_config:ocean.delta_sl.file_doc = "Name of the file containing sea level offsets.";
    pism_config:ocean.delta_sl.file_option = "ocean_delta_sl_file";
    pism_config:ocean.delta_sl.file_type = "string";

    pism_config:ocean.delta_sl.periodic = "no";
    pism_config:ocean.delta_sl.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.delta_sl.periodic_type = "flag";

    pism_config:ocean.delta_sl_2d.file = "";
    pism_config:ocean.delta_sl_2d.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:ocean.delta_sl_2d.file_type = "string";

    pism_config:ocean.delta_sl_2d.periodic = "no";
    pism_config:ocean.delta_sl_2d.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.delta_sl_2d.periodic_type = "flag";

    pism_config:ocean.frac_MBP.file = "";
    pism_config:ocean.frac_MBP.file_doc = "Name of the file containing melange back-pressure scaling.";
    pism_config:ocean.frac_MBP.file_option = "ocean_frac_MBP_file";
    pism_config:ocean.frac_MBP.file_type = "string";

    pism_config:ocean.frac_MBP.periodic = "no";
    pism_config:ocean.frac_MBP.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.frac_MBP.periodic_type = "flag";

    pism_config:ocean.frac_mass_flux.file = "";
    pism_config:ocean.frac_mass_flux.file_doc = "Name of the file containing sub-shelf mass flux scaling.";
    pism_config:ocean.frac_mass_flux.file_option = "ocean_frac_mass_flux_file";
    pism_config:ocean.frac_mass_flux.file_type = "string";

    pism_config:ocean.frac_mass_flux.periodic = "no";
    pism_config:ocean.frac_mass_flux.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.frac_mass_flux.periodic_type = "flag";

    pism_config:ocean.given.file = "";
    pism_config:ocean.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:ocean.given.file_option = "ocean_given_file";
    pism_config:ocean.given.file_type = "string";

    pism_config:ocean.given.periodic = "no";
    pism_config:ocean.given.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.given.periodic_type = "flag";

    pism_config:ocean.models = "constant";
    pism_config:ocean.models_doc = "Comma-separated list of ocean models and modifiers";
    pism_config:ocean.models_option = "ocean";
    pism_config:ocean.models_type = "string";

    pism_config:ocean.pico.continental_shelf_depth = -800.0;
    pism_config:ocean.pico.continental_shelf_depth_doc = "Specifies the depth up to which oceanic input temperatures and salinities are averaged over the continental shelf areas in front of the ice shelf cavities.";
    pism_config:ocean.pico.continental_shelf_depth_option = "continental_shelf_depth";
    pism_config:ocean.pico.continental_shelf_depth_type = "number";
    pism_config:ocean.pico.continental_shelf_depth_units = "meters";

    pism_config:ocean.pico.exclude_ice_rises = "yes";
    pism_config:ocean.pico.exclude_ice_rises_doc = "If set to true, grounding lines of ice rises are excluded in the geometrical routines that determine the ocean boxes; using this option is recommended.";
    pism_config:ocean.pico.exclude_ice_rises_option = "exclude_icerises";
    pism_config:ocean.pico.exclude_ice_rises_type = "flag";

    pism_config:ocean.pico.file = "";
    pism_config:ocean.pico.file_doc = "Specifies the NetCDF file containing potential temperature (:var:`theta_ocean`), salinity (:var:`salinity_ocean`) and ocean basins (:var:`basins`).";
    pism_config:ocean.pico.file_option = "ocean_pico_file";
    pism_config:ocean.pico.file_type = "string";

    pism_config:ocean.pico.heat_exchange_coefficent = 2e-5;
    pism_config:ocean.pico.heat_exchange_coefficent_doc = "Sets the coefficient for turbulent heat exchange from the ambient ocean across the boundary layer beneath the ice shelf base.";
    pism_config:ocean.pico.heat_exchange_coefficent_option = "gamma_T";
    pism_config:ocean.pico.heat_exchange_coefficent_type = "number";
    pism_config:ocean.pico.heat_exchange_coefficent_units = "meters second-1";

    pism_config:ocean.pico.maximum_ice_rise_area = 1e5;
    pism_config:ocean.pico.maximum_ice_rise_area_doc = "Specifies an area threshold that separates ice rises from continental regions.";
    pism_config:ocean.pico.maximum_ice_rise_area_type = "number";
    pism_config:ocean.pico.maximum_ice_rise_area_units = "km2";

    pism_config:ocean.pico.number_of_boxes = 5;
    pism_config:ocean.pico.number_of_boxes_doc = "For each ice shelf the number of ocean boxes is determined by interpolating between 1 and number_of_boxes depending on its size and geometry such that larger ice shelves are resolved with more boxes; a value of 5 is suitable for the Antarctic setup.";
    pism_config:ocean.pico.number_of_boxes_option = "number_of_boxes";
    pism_config:ocean.pico.number_of_boxes_type = "integer";
    pism_config:ocean.pico.number_of_boxes_units = "pure number";

    pism_config:ocean.pico.overturning_coefficent = 1e6;
    pism_config:ocean.pico.overturning_coefficent_doc = "Sets the overturning strength coefficient.";
    pism_config:ocean.pico.overturning_coefficent_option = "overturning_coeff";
    pism_config:ocean.pico.overturning_coefficent_type = "number";
    pism_config:ocean.pico.overturning_coefficent_units = "meters6 seconds-1 kg-1";

    pism_config:ocean.pico.periodic = "no";
    pism_config:ocean.pico.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.pico.periodic_type = "flag";

    pism_config:ocean.pik_melt_factor = 5e-3;
    pism_config:ocean.pik_melt_factor_doc = "dimensionless tuning parameter in the ``-ocean pik`` ocean heat flux parameterization; see :cite:`Martinetal2011`";
    pism_config:ocean.pik_melt_factor_option = "meltfactor_pik";
    pism_config:ocean.pik_melt_factor_type = "number";
    pism_config:ocean.pik_melt_factor_units = "1";

    pism_config:ocean.runoff_to_ocean_melt.b = 0.15;
    pism_config:ocean.runoff_to_ocean_melt.b_doc = "parameter B in eqn. 1 in :cite:`Aschwanden2019`";
    pism_config:ocean.runoff_to_ocean_melt.b_type = "number";
    pism_config:ocean.runoff_to_ocean_melt.b_units = "1";

    pism_config:ocean.runoff_to_ocean_melt.file = "";
    pism_config:ocean.runoff_to_ocean_melt.file_doc = "Name of the file containing the ``delta_T`` variable used to scale ocean melt";
    pism_config:ocean.runoff_to_ocean_melt.file_option = "ocean_runoff_smb";
    pism_config:ocean.runoff_to_ocean_melt.file_type = "string";

    pism_config:ocean.runoff_to_ocean_melt.power_alpha = 0.54;
    pism_config:ocean.runoff_to_ocean_melt.power_alpha_doc = "exponent `\\alpha` in eqn. 1 in :cite:`Xu2013`";
    pism_config:ocean.runoff_to_ocean_melt.power_alpha_type = "number";
    pism_config:ocean.runoff_to_ocean_melt.power_alpha_units = "1";

    pism_config:ocean.runoff_to_ocean_melt.power_beta = 1.17;
    pism_config:ocean.runoff_to_ocean_melt.power_beta_doc = "exponent `\\beta` in eqn. 1 in :cite:`Xu2013`";
    pism_config:ocean.runoff_to_ocean_melt.power_beta_type = "number";
    pism_config:ocean.runoff_to_ocean_melt.power_beta_units = "1";

    pism_config:ocean.sub_shelf_heat_flux_into_ice = 0.5;
    pism_config:ocean.sub_shelf_heat_flux_into_ice_doc = "= J meter-2 second-1; naively chosen default value for heat from ocean; see comments in pism::ocean::Constant::shelf_base_mass_flux().";
    pism_config:ocean.sub_shelf_heat_flux_into_ice_type = "number";
    pism_config:ocean.sub_shelf_heat_flux_into_ice_units = "W meter-2";

    pism_config:ocean.th.clip_salinity = "yes";
    pism_config:ocean.th.clip_salinity_doc = "Clip shelf base salinity so that it is in the range [4, 40] k/kg. See :cite:`HollandJenkins1999`.";
    pism_config:ocean.th.clip_salinity_option = "clip_shelf_base_salinity";
    pism_config:ocean.th.clip_salinity_type = "flag";

    pism_config:ocean.th.file = "";
    pism_config:ocean.th.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:ocean.th.file_option = "ocean_th_file";
    pism_config:ocean.th.file_type = "string";

    pism_config:ocean.th.gamma_S = 5.05e-7;
    pism_config:ocean.th.gamma_S_doc = "Turbulent salt transfer coefficient. See :cite:`HollandJenkins1999`.";
    pism_config:ocean.th.gamma_S_option = "gamma_T";
    pism_config:ocean.th.gamma_S_type = "number";
    pism_config:ocean.th.gamma_S_units = "m s-1";

    pism_config:ocean.th.gamma_T = 1.00e-4;
    pism_config:ocean.th.gamma_T_doc = "Turbulent heat transfer coefficient. See :cite:`HollandJenkins1999`.";
    pism_config:ocean.th.gamma_T_option = "gamma_T";
    pism_config:ocean.th.gamma_T_type = "number";
    pism_config:ocean.th.gamma_T_units = "m s-1";

    pism_config:ocean.th.periodic = "no";
    pism_config:ocean.th.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:ocean.th.periodic_type = "flag";

    pism_config:output.ISMIP6 = "false";
    pism_config:output.ISMIP6_doc = "Follow ISMIP6 conventions (units, variable names, \"standard names\") when writing output variables.";
    pism_config:output.ISMIP6_type = "flag";

    pism_config:output.ISMIP6_extra_variables = "lithk,orog,topg,hfgeoubed,acabf,libmassbfgr,libmassbffl,dlithkdt,velsurf,zvelsurf,velbase,zvelbase,velmean,litemptop,litempbotgr,litempbotfl,strbasemag,licalvf,lifmassbf,sftgif,sftgrf,sftflf";
    pism_config:output.ISMIP6_extra_variables_doc = "Comma-separated list of fields reported by models participating in ISMIP6 simulations.";
    pism_config:output.ISMIP6_extra_variables_type = "string";

    pism_config:output.ISMIP6_ts_variables = "lim,limnsw,iareagr,iareafl,tendacabf,tendlibmassbf,tendlibmassbffl,tendlicalvf,tendlifmassbf";
    pism_config:output.ISMIP6_ts_variables_doc = "Comma-separated list of scalar variables (time series) reported by models participating in ISMIP6 simulations.";
    pism_config:output.ISMIP6_ts_variables_type = "string";

    pism_config:output.checkpoint.exit = "no";
    pism_config:output.checkpoint.exit_doc = "If ``true`` PISM will exit with after checkpointing.";
    pism_config:output.checkpoint.exit_type = "flag";

    pism_config:output.checkpoint.exit_code = 85;
    pism_config:output.checkpoint.exit_code_doc = "Exit code to use if :config:`output.checkpoint.exit` is set.";
    pism_config:output.checkpoint.exit_code_type = "integer";
    pism_config:output.checkpoint.exit_code_units = "none";

    pism_config:output.checkpoint.file = "";
    pism_config:output.checkpoint.file_doc = "If set, save model checkpoints to this file, otherwise build the name by appending ``_checkpoint`` to :config:`output.file`.";
    pism_config:output.checkpoint.file_type = "string";

    pism_config:output.checkpoint.interval = 1.0;
    pism_config:output.checkpoint.interval_doc = "wall-clock time between checkpointing";
    pism_config:output.checkpoint.interval_option = "checkpoint_interval";
    pism_config:output.checkpoint.interval_type = "number";
    pism_config:output.checkpoint.interval_units = "hours";

    pism_config:output.checkpoint.size = "small";
    pism_config:output.checkpoint.size_choices = "none,small,medium,big_2d,big";
    pism_config:output.checkpoint.size_doc = "The \"size\" of a checkpoint file. See parameters :config:`output.sizes.medium`, :config:`output.sizes.big_2d`, :config:`output.sizes.big`";
    pism_config:output.checkpoint.size_option = "checkpoint_size";
    pism_config:output.checkpoint.size_type = "keyword";

    pism_config:output.compression_level = 0;
    pism_config:output.compression_level_doc = "Compression level for 2D and 3D output variables (if supported by :config:`output.format`)";
    pism_config:output.compression_level_type = "integer";
    pism_config:output.compression_level_units = "count";

    pism_config:output.extra.append = "no";
    pism_config:output.extra.append_doc = "Append to an existing output file.  No effect if file does not yet exist, and no effect if :config:`output.extra.split` is set.";
    pism_config:output.extra.append_option = "extra_append";
    pism_config:output.extra.append_type = "flag";

    pism_config:output.extra.file = "";
    pism_config:output.extra.file_doc = "Name of the file that will contain spatially-variable diagnostics. Should be different from :config:`output.file`.";
    pism_config:output.extra.file_option = "extra_file";
    pism_config:output.extra.file_type = "string";

    pism_config:output.extra.split = "no";
    pism_config:output.extra.split_doc = "Save spatially-variable diagnostics to separate files (one per time record).";
    pism_config:output.extra.split_option = "extra_split";
    pism_config:output.extra.split_type = "flag";

    pism_config:output.extra.stop_missing = "yes";
    pism_config:output.extra.stop_missing_doc = "Stop if requested variable is not available instead of warning.";
    pism_config:output.extra.stop_missing_option = "extra_stop_missing";
    pism_config:output.extra.stop_missing_type = "flag";

    pism_config:output.extra.times = "";
    pism_config:output.extra.times_doc = "List or a range of times defining reporting intervals for spatially-variable diagnostics.";
    pism_config:output.extra.times_option = "extra_times";
    pism_config:output.extra.times_type = "string";

    pism_config:output.extra.vars = "";
    pism_config:output.extra.vars_doc = "Comma-separated list of spatially-variable diagnostics.";
    pism_config:output.extra.vars_option = "extra_vars";
    pism_config:output.extra.vars_type = "string";

    pism_config:output.file = "unnamed.nc";
    pism_config:output.file_doc = "The file to save final model results to.";
    pism_config:output.file_option = "o";
    pism_config:output.file_type = "string";

    pism_config:output.fill_value = -2e9;
    pism_config:output.fill_value_doc = "_FillValue used when saving diagnostic quantities";
    pism_config:output.fill_value_type = "number";
    pism_config:output.fill_value_units = "none";

    pism_config:output.format = "netcdf3";
    pism_config:output.format_choices = "netcdf3,netcdf4_serial,netcdf4_parallel,pnetcdf,pio_pnetcdf,pio_netcdf4p,pio_netcdf4c,pio_netcdf";
    pism_config:output.format_doc = "The I/O format used for spatial fields; ``netcdf3`` is the default, ``netcd4_parallel`` is available if PISM was built with parallel NetCDF-4, and ``pnetcdf`` is available if PISM was built with PnetCDF.";
    pism_config:output.format_option = "o_format";
    pism_config:output.format_type = "keyword";

    pism_config:output.ice_free_thickness_standard = 10.0;
    pism_config:output.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a grid cell is considered ice-free for purposes of reporting glacierized area, volume, etc.";
    pism_config:output.ice_free_thickness_standard_type = "number";
    pism_config:output.ice_free_thickness_standard_units = "meters";

    pism_config:output.pio.base = 0;
    pism_config:output.pio.base_doc = "Rank of the first I/O task";
    pism_config:output.pio.base_type = "integer";
    pism_config:output.pio.base_units = "count";

    pism_config:output.pio.n_writers = 1;
    pism_config:output.pio.n_writers_doc = "Number of I/O tasks to use";
    pism_config:output.pio.n_writers_type = "integer";
    pism_config:output.pio.n_writers_units = "count";

    pism_config:output.pio.stride = 1;
    pism_config:output.pio.stride_doc = "Offset between I/O tasks";
    pism_config:output.pio.stride_type = "integer";
    pism_config:output.pio.stride_units = "count";

    pism_config:output.runtime.area_scale_factor_log10 = 6;
    pism_config:output.runtime.area_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for area (in km^2) in summary line to stdout";
    pism_config:output.runtime.area_scale_factor_log10_option = "summary_area_scale_factor_log10";
    pism_config:output.runtime.area_scale_factor_log10_type = "integer";
    pism_config:output.runtime.area_scale_factor_log10_units = "pure number";

    pism_config:output.runtime.time_unit_name = "year";
    pism_config:output.runtime.time_unit_name_doc = "Time units used when printing model time, time step, and maximum horizontal velocity at summary to stdout.  Must be valid udunits for time.  (E.g. choose from year,month,day,hour,minute,second.)";
    pism_config:output.runtime.time_unit_name_type = "string";

    pism_config:output.runtime.time_use_calendar = "yes";
    pism_config:output.runtime.time_use_calendar_doc = "Whether to use the current calendar when printing model time in summary to stdout.";
    pism_config:output.runtime.time_use_calendar_type = "flag";

    pism_config:output.runtime.viewer.size = 320;
    pism_config:output.runtime.viewer.size_doc = "default diagnostic viewer size (number of pixels of the longer side)";
    pism_config:output.runtime.viewer.size_option = "view_size";
    pism_config:output.runtime.viewer.size_type = "integer";
    pism_config:output.runtime.viewer.size_units = "count";

    pism_config:output.runtime.viewer.variables = "";
    pism_config:output.runtime.viewer.variables_doc = "comma-separated list of map-plane diagnostic quantities to view at runtime";
    pism_config:output.runtime.viewer.variables_option = "view";
    pism_config:output.runtime.viewer.variables_type = "string";

    pism_config:output.runtime.volume_scale_factor_log10 = 6;
    pism_config:output.runtime.volume_scale_factor_log10_doc = "an integer; log base 10 of scale factor to use for volume (in km^3) in summary line to stdout";
    pism_config:output.runtime.volume_scale_factor_log10_option = "summary_vol_scale_factor_log10";
    pism_config:output.runtime.volume_scale_factor_log10_type = "integer";
    pism_config:output.runtime.volume_scale_factor_log10_units = "pure number";

    pism_config:output.size = "medium";
    pism_config:output.size_choices = "none,small,medium,big_2d,big";
    pism_config:output.size_doc = "The \"size\" of an output file. See parameters :config:`output.sizes.medium`, :config:`output.sizes.big_2d`, :config:`output.sizes.big`";
    pism_config:output.size_option = "o_size";
    pism_config:output.size_type = "keyword";

    pism_config:output.sizes.big = "cts,liqfrac,temp,temp_pa,uvel,vvel,wvel,wvel_rel";
    pism_config:output.sizes.big_doc = "Comma-separated list of variables to write to the output (in addition to ``model_state`` variables and variables listed in :config:`output.sizes.medium` and :config:`output.sizes.big_2d`) if ``big`` output size is selected. Does not include fields written by sub-models.";
    pism_config:output.sizes.big_type = "string";

    pism_config:output.sizes.big_2d = "age,bfrict,bheatflx,bmelt,bwp,bwprel,dbdt,effbwp,enthalpybase,enthalpysurf,flux_divergence,hardav,hydroinput,lat,litho_temp,lon,nuH,rank,tempbase,tempicethk,tempicethk_basal,temppabase,tempsurf,thk,thksmooth,tillphi,topg,velbar,velbase,wallmelt,wvelbase";
    pism_config:output.sizes.big_2d_doc = "Comma-separated list of variables to write to the output (in addition to ``model_state`` variables and variables listed in :config:`output.sizes.medium`) if ``big_2d`` output size is selected. Does not include fields written by boundary models.";
    pism_config:output.sizes.big_2d_type = "string";

    pism_config:output.sizes.medium = "bwat,bwatvel,climatic_mass_balance,diffusivity,enthalpy,flux,flux_mag,ice_surface_temp,liqfrac,mask,schoofs_theta,strain_rates,taub_mag,tauc,taud_mag,temp_pa,tillwat,topgsmooth,usurf,velbar_mag,velbase_mag,velsurf,velsurf_mag,wvelsurf";
    pism_config:output.sizes.medium_doc = "Comma-separated list of variables to write to the output (in addition to ``model_state`` variables) if ``medium`` output size (the default) is selected. Does not include fields written by sub-models.";
    pism_config:output.sizes.medium_type = "string";

    pism_config:output.snapshot.file = "";
    pism_config:output.snapshot.file_doc = "Snapshot (output) file name (or prefix, if saving to individual files).";
    pism_config:output.snapshot.file_option = "save_file";
    pism_config:output.snapshot.file_type = "string";

    pism_config:output.snapshot.size = "small";
    pism_config:output.snapshot.size_choices = "none,small,medium,big_2d,big";
    pism_config:output.snapshot.size_doc = "The \"size\" of a snapshot file. See parameters :config:`output.sizes.medium`, :config:`output.sizes.big_2d`, :config:`output.sizes.big`";
    pism_config:output.snapshot.size_option = "save_size";
    pism_config:output.snapshot.size_type = "keyword";

    pism_config:output.snapshot.split = "no";
    pism_config:output.snapshot.split_doc = "Save model state snapshots to separate files (one per time record).";
    pism_config:output.snapshot.split_option = "save_split";
    pism_config:output.snapshot.split_type = "flag";

    pism_config:output.snapshot.times = "";
    pism_config:output.snapshot.times_doc = "List or a range of times to save model state snapshots at.";
    pism_config:output.snapshot.times_option = "save_times";
    pism_config:output.snapshot.times_type = "string";

    pism_config:output.timeseries.append = "false";
    pism_config:output.timeseries.append_doc = "If true, append to the scalar time series output file.";
    pism_config:output.timeseries.append_option = "ts_append";
    pism_config:output.timeseries.append_type = "flag";

    pism_config:output.timeseries.buffer_size = 10000;
    pism_config:output.timeseries.buffer_size_doc = "Number of scalar diagnostic time-series records to hold in memory before writing to disk. (PISM writes this many time-series records to reduce I/O costs.) Send the USR2 signal to flush time-series.";
    pism_config:output.timeseries.buffer_size_type = "integer";
    pism_config:output.timeseries.buffer_size_units = "count";

    pism_config:output.timeseries.filename = "";
    pism_config:output.timeseries.filename_doc = "Name of the file to save scalar time series to. Leave empty to disable reporting scalar time-series.";
    pism_config:output.timeseries.filename_option = "ts_file";
    pism_config:output.timeseries.filename_type = "string";

    pism_config:output.timeseries.times = "";
    pism_config:output.timeseries.times_doc = "List or range of times defining reporting time intervals.";
    pism_config:output.timeseries.times_option = "ts_times";
    pism_config:output.timeseries.times_type = "string";

    pism_config:output.timeseries.variables = "";
    pism_config:output.timeseries.variables_doc = "Requested scalar (time-series) diagnostics. Leave empty to save all available diagnostics.";
    pism_config:output.timeseries.variables_option = "ts_vars";
    pism_config:output.timeseries.variables_type = "string";

    pism_config:output.use_MKS = "false";
    pism_config:output.use_MKS_doc = "Use MKS units in output files.";
    pism_config:output.use_MKS_type = "flag";

    pism_config:regional.no_model_strip = 5.0;
    pism_config:regional.no_model_strip_doc = "Default width of the \"no model strip\" in regional setups.";
    pism_config:regional.no_model_strip_option = "no_model_strip";
    pism_config:regional.no_model_strip_type = "number";
    pism_config:regional.no_model_strip_units = "km";

    pism_config:regional.no_model_yield_stress = 1000.0;
    pism_config:regional.no_model_yield_stress_doc = "High yield stress used in the ``no_model_mask`` area in the regional mode.";
    pism_config:regional.no_model_yield_stress_type = "number";
    pism_config:regional.no_model_yield_stress_units = "kPa";

    pism_config:regional.zero_gradient = "false";
    pism_config:regional.zero_gradient_doc = "Use zero ice thickness and ice surface gradient in the no_model_mask area.";
    pism_config:regional.zero_gradient_option = "zero_grad_where_no_model";
    pism_config:regional.zero_gradient_type = "flag";

    pism_config:run_info.institution = "";
    pism_config:run_info.institution_doc = "Institution name. This string is written to output files as the ``institution`` global attribute.";
    pism_config:run_info.institution_option = "institution";
    pism_config:run_info.institution_type = "string";

    pism_config:run_info.title = "";
    pism_config:run_info.title_doc = "Free-form string containing a concise description of the current run. This string is written to output files as the ``title`` global attribute.";
    pism_config:run_info.title_option = "title";
    pism_config:run_info.title_type = "string";

    pism_config:sea_level.constant.value = 0.0;
    pism_config:sea_level.constant.value_doc = "Sea level elevation used by the ``constant`` sea level model";
    pism_config:sea_level.constant.value_units = "meters";
    pism_config:sea_level.constant.value_type = "number";

    pism_config:sea_level.models = "constant";
    pism_config:sea_level.models_doc = "Comma-separated list of sea level models and modifiers";
    pism_config:sea_level.models_option = "sea_level";
    pism_config:sea_level.models_type = "string";

    pism_config:stress_balance.blatter.Glen_exponent_units = "pure number";
    pism_config:stress_balance.blatter.Glen_exponent_type = "number";
    pism_config:stress_balance.blatter.Glen_exponent = 3.0;
    pism_config:stress_balance.blatter.Glen_exponent_doc = "Glen exponent in ice flow law for the Blatter stress balance solver";

    pism_config:stress_balance.blatter.Mz_option = "blatter_Mz";
    pism_config:stress_balance.blatter.Mz_units = "count";
    pism_config:stress_balance.blatter.Mz_type = "integer";
    pism_config:stress_balance.blatter.Mz = 5;
    pism_config:stress_balance.blatter.Mz_doc = "Number of vertical grid levels in the ice";

    pism_config:stress_balance.blatter.coarsening_factor_option = "blatter_coarsening_factor";
    pism_config:stress_balance.blatter.coarsening_factor_units = "count";
    pism_config:stress_balance.blatter.coarsening_factor_type = "integer";
    pism_config:stress_balance.blatter.coarsening_factor = 2;
    pism_config:stress_balance.blatter.coarsening_factor_doc = "Coarsening factor in the `z` direction";

    pism_config:stress_balance.blatter.enhancement_factor_option = "blatter_e";
    pism_config:stress_balance.blatter.enhancement_factor_units = "1";
    pism_config:stress_balance.blatter.enhancement_factor_type = "number";
    pism_config:stress_balance.blatter.enhancement_factor = 1.0;
    pism_config:stress_balance.blatter.enhancement_factor_doc = "Flow enhancement factor for the Blatter stress balance flow law";

    pism_config:stress_balance.blatter.flow_law_type = "keyword";
    pism_config:stress_balance.blatter.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb";
    pism_config:stress_balance.blatter.flow_law = "gpbld";
    pism_config:stress_balance.blatter.flow_law_doc = "The flow law used by the Blatter-Pattyn stress balance model";

    pism_config:stress_balance.blatter.use_eta_transform_type = "flag";
    pism_config:stress_balance.blatter.use_eta_transform = "no";
    pism_config:stress_balance.blatter.use_eta_transform_doc = "Use the `\\eta` transform to improve the accuracy of the surface gradient approximation near grounded margins (see :cite:`BLKCB` for details).";

    pism_config:stress_balance.calving_front_stress_bc = "no";
    pism_config:stress_balance.calving_front_stress_bc_doc = "Apply CFBC condition as in :cite:`Albrechtetal2011`, :cite:`Winkelmannetal2011`.  May only apply to some stress balances; e.g. SSAFD as of May 2011.  If not set then a strength-extension is used, as in :cite:`BBssasliding`.";
    pism_config:stress_balance.calving_front_stress_bc_option = "cfbc";
    pism_config:stress_balance.calving_front_stress_bc_type = "flag";

    pism_config:stress_balance.ice_free_thickness_standard = 10.0;
    pism_config:stress_balance.ice_free_thickness_standard_doc = "If ice is thinner than this standard then a cell is considered ice-free for purposes of computing ice velocity distribution.";
    pism_config:stress_balance.ice_free_thickness_standard_type = "number";
    pism_config:stress_balance.ice_free_thickness_standard_units = "meters";

    pism_config:stress_balance.model = "sia";
    pism_config:stress_balance.model_choices = "none,prescribed_sliding,weertman_sliding,sia,ssa,prescribed_sliding+sia,weertman_sliding+sia,ssa+sia,blatter";
    pism_config:stress_balance.model_doc = "Stress balance model";
    pism_config:stress_balance.model_option = "stress_balance";
    pism_config:stress_balance.model_type = "keyword";

    pism_config:stress_balance.prescribed_sliding.file = "";
    pism_config:stress_balance.prescribed_sliding.file_doc = "The name of the file containing prescribed sliding velocity (variable names: :var:`ubar`, :var:`vbar`).";
    pism_config:stress_balance.prescribed_sliding.file_type = "string";

    pism_config:stress_balance.sia.Glen_exponent = 3.0;
    pism_config:stress_balance.sia.Glen_exponent_doc = "Glen exponent in ice flow law for SIA";
    pism_config:stress_balance.sia.Glen_exponent_option = "sia_n";
    pism_config:stress_balance.sia.Glen_exponent_type = "number";
    pism_config:stress_balance.sia.Glen_exponent_units = "pure number";

    pism_config:stress_balance.sia.bed_smoother.range = 5.0e3;
    pism_config:stress_balance.sia.bed_smoother.range_doc = "half-width of smoothing domain in the bed roughness parameterization for SIA :cite:`Schoofbasaltopg2003`; set to zero to disable";
    pism_config:stress_balance.sia.bed_smoother.range_option = "bed_smoother_range";
    pism_config:stress_balance.sia.bed_smoother.range_type = "number";
    pism_config:stress_balance.sia.bed_smoother.range_units = "meters";

    pism_config:stress_balance.sia.bed_smoother.theta_min = 0.0;
    pism_config:stress_balance.sia.bed_smoother.theta_min_doc = "minimum value of `\\theta` in the bed roughness parameterization for SIA :cite:`Schoofbasaltopg2003`";
    pism_config:stress_balance.sia.bed_smoother.theta_min_type = "number";
    pism_config:stress_balance.sia.bed_smoother.theta_min_units = "1";

    pism_config:stress_balance.sia.e_age_coupling = "no";
    pism_config:stress_balance.sia.e_age_coupling_doc = "Couple the SIA enhancement factor to age as in :cite:`Greve`.";
    pism_config:stress_balance.sia.e_age_coupling_option = "e_age_coupling";
    pism_config:stress_balance.sia.e_age_coupling_type = "flag";

    pism_config:stress_balance.sia.enhancement_factor = 1.0;
    pism_config:stress_balance.sia.enhancement_factor_doc = "Flow enhancement factor for SIA";
    pism_config:stress_balance.sia.enhancement_factor_option = "sia_e";
    pism_config:stress_balance.sia.enhancement_factor_type = "number";
    pism_config:stress_balance.sia.enhancement_factor_units = "1";

    pism_config:stress_balance.sia.enhancement_factor_interglacial = 1.0;
    pism_config:stress_balance.sia.enhancement_factor_interglacial_doc = "Flow enhancement factor for SIA; used for ice accumulated during interglacial periods.";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_option = "sia_e_interglacial";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_type = "number";
    pism_config:stress_balance.sia.enhancement_factor_interglacial_units = "1";

    pism_config:stress_balance.sia.flow_law = "gpbld";
    pism_config:stress_balance.sia.flow_law_choices = "arr,arrwarm,gk,gpbld,hooke,isothermal_glen,pb";
    pism_config:stress_balance.sia.flow_law_doc = "The SIA flow law.";
    pism_config:stress_balance.sia.flow_law_option = "sia_flow_law";
    pism_config:stress_balance.sia.flow_law_type = "keyword";

    pism_config:stress_balance.sia.grain_size_age_coupling = "no";
    pism_config:stress_balance.sia.grain_size_age_coupling_doc = "Use age of the ice to compute grain size to use with the Goldsby-Kohlstedt :cite:`GoldsbyKohlstedt` flow law";
    pism_config:stress_balance.sia.grain_size_age_coupling_option = "grain_size_age_coupling";
    pism_config:stress_balance.sia.grain_size_age_coupling_type = "flag";

    pism_config:stress_balance.sia.limit_diffusivity = "no";
    pism_config:stress_balance.sia.limit_diffusivity_doc = "Limit SIA diffusivity by :config:`stress_balance.sia.max_diffusivity`.";
    pism_config:stress_balance.sia.limit_diffusivity_option = "limit_sia_diffusivity";
    pism_config:stress_balance.sia.limit_diffusivity_type = "flag";

    pism_config:stress_balance.sia.max_diffusivity = 100.0;
    pism_config:stress_balance.sia.max_diffusivity_doc = "Maximum allowed diffusivity of the SIA flow. PISM stops with an error message if the SIA diffusivity exceeds this limit.";
    pism_config:stress_balance.sia.max_diffusivity_type = "number";
    pism_config:stress_balance.sia.max_diffusivity_units = "m2 s-1";

    pism_config:stress_balance.sia.surface_gradient_method = "haseloff";
    pism_config:stress_balance.sia.surface_gradient_method_choices = "eta,haseloff,mahaffy";
    pism_config:stress_balance.sia.surface_gradient_method_doc = "method used for surface gradient calculation at staggered grid points";
    pism_config:stress_balance.sia.surface_gradient_method_option = "gradient";
    pism_config:stress_balance.sia.surface_gradient_method_type = "keyword";

    pism_config:stress_balance.ssa.Glen_exponent = 3.0;
    pism_config:stress_balance.ssa.Glen_exponent_doc = "Glen exponent in ice flow law for SSA";
    pism_config:stress_balance.ssa.Glen_exponent_option = "ssa_n";
    pism_config:stress_balance.ssa.Glen_exponent_type = "number";
    pism_config:stress_balance.ssa.Glen_exponent_units = "pure number";

    pism_config:stress_balance.ssa.compute_surface_gradient_inward = "no";
    pism_config:stress_balance.ssa.compute_surface_gradient_inward_doc = "If yes then use inward first-order differencing in computing surface gradient in the SSA objects.";
    pism_config:stress_balance.ssa.compute_surface_gradient_inward_type = "flag";

    pism_config:stress_balance.ssa.dirichlet_bc = "no";
    pism_config:stress_balance.ssa.dirichlet_bc_doc = "apply SSA velocity Dirichlet boundary condition";
    pism_config:stress_balance.ssa.dirichlet_bc_option = "ssa_dirichlet_bc";
    pism_config:stress_balance.ssa.dirichlet_bc_type = "flag";

    pism_config:stress_balance.ssa.enhancement_factor = 1.0;
    pism_config:stress_balance.ssa.enhancement_factor_doc = "Flow enhancement factor for SSA";
    pism_config:stress_balance.ssa.enhancement_factor_option = "ssa_e";
    pism_config:stress_balance.ssa.enhancement_factor_type = "number";
    pism_config:stress_balance.ssa.enhancement_factor_units = "1";

    pism_config:stress_balance.ssa.epsilon = 1.0e13;
    pism_config:stress_balance.ssa.epsilon_doc = "Initial amount of regularization in computation of product of effective viscosity and thickness (`\\nu H`).  This default value for `\\nu H` comes e.g. from a hardness for the Ross ice shelf (`\\bar B`) = 1.9e8 Pa `s^{1/3}` :cite:`MacAyealetal` and a typical strain rate of 0.001 1/year for the Ross ice shelf, giving `\\nu = (\\bar B) / (2 \\cdot 0.001^{2/3})` = 9.49e+14 Pa s ~ 30 MPa year, the value in :cite:`Ritzetal2001`, but with a tiny thickness `H` of about 1 cm.";
    pism_config:stress_balance.ssa.epsilon_option = "ssa_eps";
    pism_config:stress_balance.ssa.epsilon_type = "number";
    pism_config:stress_balance.ssa.epsilon_units = "Pascal second meter";

    pism_config:stress_balance.ssa.fd.absolute_tolerance = 100.0;
    pism_config:stress_balance.ssa.fd.absolute_tolerance_doc = "Absolute tolerance used by the SNES-based SSAFD solver (converged if the infinity norm of the residual is below this)";
    pism_config:stress_balance.ssa.fd.absolute_tolerance_type = "number";
    pism_config:stress_balance.ssa.fd.absolute_tolerance_units = "Pascal";

    pism_config:stress_balance.ssa.fd.brutal_sliding = "false";
    pism_config:stress_balance.ssa.fd.brutal_sliding_doc = "Enhance sliding speed brutally.";
    pism_config:stress_balance.ssa.fd.brutal_sliding_option = "brutal_sliding";
    pism_config:stress_balance.ssa.fd.brutal_sliding_type = "flag";

    pism_config:stress_balance.ssa.fd.brutal_sliding_scale = 1.0;
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_doc = "Brutal SSA Sliding Scale";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_option = "brutal_sliding_scale";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_type = "number";
    pism_config:stress_balance.ssa.fd.brutal_sliding_scale_units = "1";

    pism_config:stress_balance.ssa.fd.extrapolate_at_margins = "true";
    pism_config:stress_balance.ssa.fd.extrapolate_at_margins_doc = "Extrapolate SSA velocity to ice-free cells near the margin to improve SSA velocities at advancing ice fronts";
    pism_config:stress_balance.ssa.fd.extrapolate_at_margins_type = "flag";

    pism_config:stress_balance.ssa.fd.flow_line_mode = "false";
    pism_config:stress_balance.ssa.fd.flow_line_mode_doc = "Set `v` (the `y` component of the ice velocity) to zero when assembling the system";
    pism_config:stress_balance.ssa.fd.flow_line_mode_type = "flag";

    pism_config:stress_balance.ssa.fd.lateral_drag.enabled = "false";
    pism_config:stress_balance.ssa.fd.lateral_drag.enabled_doc = "Set viscosity at ice shelf margin next to ice free bedrock as friction parameterization";
    pism_config:stress_balance.ssa.fd.lateral_drag.enabled_type = "flag";

    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity = 5.0e15;
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_doc = "Staggered viscosity used as side friction parameterization.";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_option = "nu_bedrock";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_type = "number";
    pism_config:stress_balance.ssa.fd.lateral_drag.viscosity_units = "Pascal second";

    pism_config:stress_balance.ssa.fd.max_iterations = 300;
    pism_config:stress_balance.ssa.fd.max_iterations_doc = "Maximum number of Picard iterations for the ice viscosity computation, in the ``SSAFD`` object";
    pism_config:stress_balance.ssa.fd.max_iterations_option = "ssafd_picard_maxi";
    pism_config:stress_balance.ssa.fd.max_iterations_type = "integer";
    pism_config:stress_balance.ssa.fd.max_iterations_units = "count";

    pism_config:stress_balance.ssa.fd.max_speed = 300000;
    pism_config:stress_balance.ssa.fd.max_speed_doc = "Upper bound for the ice speed computed by the ``SSAFD`` solver.";
    pism_config:stress_balance.ssa.fd.max_speed_option = "ssafd_max_speed";
    pism_config:stress_balance.ssa.fd.max_speed_type = "number";
    pism_config:stress_balance.ssa.fd.max_speed_units = "km s-1";

    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation = 0.8;
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_doc = "In event of \"Effective viscosity not converged\" failure, use outer iteration rule nuH <- nuH + f (nuH - nuH_old), where f is this parameter.";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_option = "ssafd_nuH_iter_failure_underrelaxation";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_type = "number";
    pism_config:stress_balance.ssa.fd.nuH_iter_failure_underrelaxation_units = "pure number";

    pism_config:stress_balance.ssa.fd.relative_convergence = 1.0e-4;
    pism_config:stress_balance.ssa.fd.relative_convergence_doc = "Relative change tolerance for the effective viscosity in the ``SSAFD`` object";
    pism_config:stress_balance.ssa.fd.relative_convergence_option = "ssafd_picard_rtol";
    pism_config:stress_balance.ssa.fd.relative_convergence_type = "number";
    pism_config:stress_balance.ssa.fd.relative_convergence_units = "1";

    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries = "yes";
    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries_doc = "Replace zero diagonal entries in the ``SSAFD`` matrix with :config:'basal_resistance.beta_ice_free_bedrock' to avoid solver failures.";
    pism_config:stress_balance.ssa.fd.replace_zero_diagonal_entries_type = "flag";

    pism_config:stress_balance.ssa.flow_law = "gpbld";
    pism_config:stress_balance.ssa.flow_law_choices = "arr,arrwarm,gpbld,hooke,isothermal_glen,pb";
    pism_config:stress_balance.ssa.flow_law_doc = "The SSA flow law.";
    pism_config:stress_balance.ssa.flow_law_option = "ssa_flow_law";
    pism_config:stress_balance.ssa.flow_law_type = "keyword";

    pism_config:stress_balance.ssa.method = "fd";
    pism_config:stress_balance.ssa.method_choices = "fd,fd_snes,fem";
    pism_config:stress_balance.ssa.method_doc = "Algorithm for computing the SSA solution.";
    pism_config:stress_balance.ssa.method_option = "ssa_method";
    pism_config:stress_balance.ssa.method_type = "keyword";

    pism_config:stress_balance.ssa.read_initial_guess = "yes";
    pism_config:stress_balance.ssa.read_initial_guess_doc = "Read the initial guess from the input file when re-starting.";
    pism_config:stress_balance.ssa.read_initial_guess_option = "ssa_read_initial_guess";
    pism_config:stress_balance.ssa.read_initial_guess_type = "flag";

    pism_config:stress_balance.ssa.strength_extension.constant_nu = 9.48680701906572e+14;
    pism_config:stress_balance.ssa.strength_extension.constant_nu_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  This value for nu comes from hardness (bar B)=1.9e8 `Pa s^{1/3}` :cite:`MacAyealetal` and a typical strain rate of 0.001 year-1:  `\\nu = (\\bar B) / (2 \\cdot 0.001^{2/3})`.  Compare the value of 9.45e14 Pa s = 30 MPa year in :cite:`Ritzetal2001`.";
    pism_config:stress_balance.ssa.strength_extension.constant_nu_type = "number";
    pism_config:stress_balance.ssa.strength_extension.constant_nu_units = "Pascal second";

    pism_config:stress_balance.ssa.strength_extension.min_thickness = 50.0;
    pism_config:stress_balance.ssa.strength_extension.min_thickness_doc = "The SSA is made elliptic by use of a constant value for the product of viscosity (nu) and thickness (H).  At ice thicknesses below this value the product nu*H switches from the normal vertical integral to a constant value.  The geometry itself is not affected by this value.";
    pism_config:stress_balance.ssa.strength_extension.min_thickness_type = "number";
    pism_config:stress_balance.ssa.strength_extension.min_thickness_units = "meters";

    pism_config:stress_balance.vertical_velocity_approximation = "centered";
    pism_config:stress_balance.vertical_velocity_approximation_choices = "centered,upstream";
    pism_config:stress_balance.vertical_velocity_approximation_doc = "Vertical velocity FD approximation. \"Upstream\" uses first-order finite difference to compute u_x and v_y. Uses basal velocity to make decisions.";
    pism_config:stress_balance.vertical_velocity_approximation_option = "vertical_velocity_approximation";
    pism_config:stress_balance.vertical_velocity_approximation_type = "keyword";

    pism_config:stress_balance.weertman_sliding.A = 1.8e-16;
    pism_config:stress_balance.weertman_sliding.A_doc = "Sliding parameter in the Weertman-style sliding parameterization :cite:`Tomkin2007`";
    pism_config:stress_balance.weertman_sliding.A_type = "number";
    pism_config:stress_balance.weertman_sliding.A_units = "Pa-3 year-1 m-2";

    pism_config:stress_balance.weertman_sliding.k = 0.2;
    pism_config:stress_balance.weertman_sliding.k_doc = "The ratio of the basal water pressure and the ice overburden pressure in the Weertman-style sliding parameterization.";
    pism_config:stress_balance.weertman_sliding.k_type = "number";
    pism_config:stress_balance.weertman_sliding.k_units = "1";

    pism_config:surface.anomaly.file = "";
    pism_config:surface.anomaly.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:surface.anomaly.file_option = "surface_anomaly_file";
    pism_config:surface.anomaly.file_type = "string";

    pism_config:surface.anomaly.periodic = "no";
    pism_config:surface.anomaly.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.anomaly.periodic_type = "flag";

    pism_config:surface.cache.update_interval = 10;
    pism_config:surface.cache.update_interval_doc = "Update interval (in 365-day years) for the ``-surface cache`` modifier.";
    pism_config:surface.cache.update_interval_type = "integer";
    pism_config:surface.cache.update_interval_units = "365days";

    pism_config:surface.debm_simple.air_temp_all_precip_as_rain = 275.15;
    pism_config:surface.debm_simple.air_temp_all_precip_as_rain_doc = "Threshold temperature above which all precipitation is interpreted as rain; must exceed :config:`surface.debm_simple.air_temp_all_precip_as_snow`";
    pism_config:surface.debm_simple.air_temp_all_precip_as_rain_type = "number";
    pism_config:surface.debm_simple.air_temp_all_precip_as_rain_units = "Kelvin";

    pism_config:surface.debm_simple.air_temp_all_precip_as_snow = 273.15;
    pism_config:surface.debm_simple.air_temp_all_precip_as_snow_doc = "Threshold temperature below which all precipitation is interpreted as snow";
    pism_config:surface.debm_simple.air_temp_all_precip_as_snow_type = "number";
    pism_config:surface.debm_simple.air_temp_all_precip_as_snow_units = "Kelvin";

    pism_config:surface.debm_simple.albedo_input.file = "";
    pism_config:surface.debm_simple.albedo_input.file_doc = "Name of the file containing the variable :var:`albedo` to use instead of parameterizing it";
    pism_config:surface.debm_simple.albedo_input.file_type = "string";

    pism_config:surface.debm_simple.albedo_input.periodic = "no";
    pism_config:surface.debm_simple.albedo_input.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.debm_simple.albedo_input.periodic_type = "flag";

    pism_config:surface.debm_simple.albedo_max = 0.82;
    pism_config:surface.debm_simple.albedo_max_doc = "Maximum (\"fresh snow\") albedo in albedo parametrization (tuning parameter)";
    pism_config:surface.debm_simple.albedo_max_type = "number";
    pism_config:surface.debm_simple.albedo_max_units = "1";

    pism_config:surface.debm_simple.albedo_min = 0.47;
    pism_config:surface.debm_simple.albedo_min_doc = "Minimum (\"bare ice\") albedo in albedo parametrization";
    pism_config:surface.debm_simple.albedo_min_type = "number";
    pism_config:surface.debm_simple.albedo_min_units = "1";

    pism_config:surface.debm_simple.albedo_ocean = 0.1;
    pism_config:surface.debm_simple.albedo_ocean_doc = "Albedo of ice-free ocean";
    pism_config:surface.debm_simple.albedo_ocean_type = "number";
    pism_config:surface.debm_simple.albedo_ocean_units = "1";

    pism_config:surface.debm_simple.albedo_slope = -790;
    pism_config:surface.debm_simple.albedo_slope_doc = "Slope in albedo parametrization (tuning parameter)";
    pism_config:surface.debm_simple.albedo_slope_type = "number";
    pism_config:surface.debm_simple.albedo_slope_units = "m2 s kg-1";

    pism_config:surface.debm_simple.c1 = 29.0;
    pism_config:surface.debm_simple.c1_doc = "Tuning parameter in the temperature-driven melt contribution";
    pism_config:surface.debm_simple.c1_type = "number";
    pism_config:surface.debm_simple.c1_units = "W m-2 K-1";

    pism_config:surface.debm_simple.c2 = -93.0;
    pism_config:surface.debm_simple.c2_doc = "Tuning parameter controlling the melt offset";
    pism_config:surface.debm_simple.c2_type = "number";
    pism_config:surface.debm_simple.c2_units = "W m-2";

    pism_config:surface.debm_simple.interpret_precip_as_snow = "no";
    pism_config:surface.debm_simple.interpret_precip_as_snow_doc = "If true, interpret *all* precipitation as snow";
    pism_config:surface.debm_simple.interpret_precip_as_snow_type = "flag";

    pism_config:surface.debm_simple.max_evals_per_year = 52;
    pism_config:surface.debm_simple.max_evals_per_year_doc = "Maximum number of air temperature and precipitation samples per year used to build location-dependent time series for computing melt and snow accumulation; the default means use weekly samples of the annual cycle";
    pism_config:surface.debm_simple.max_evals_per_year_type = "integer";
    pism_config:surface.debm_simple.max_evals_per_year_units = "count";

    pism_config:surface.debm_simple.melting_threshold_temp = 266.65;
    pism_config:surface.debm_simple.melting_threshold_temp_doc = "Threshold temperature below which no melting occurs";
    pism_config:surface.debm_simple.melting_threshold_temp_type = "number";
    pism_config:surface.debm_simple.melting_threshold_temp_units = "Kelvin";

    pism_config:surface.debm_simple.paleo.eccentricity =  0.0167;
    pism_config:surface.debm_simple.paleo.eccentricity_doc = "Eccentricity of the Earth's orbit";
    pism_config:surface.debm_simple.paleo.eccentricity_type = "number";
    pism_config:surface.debm_simple.paleo.eccentricity_units = "1";

    pism_config:surface.debm_simple.paleo.enabled = "false";
    pism_config:surface.debm_simple.paleo.enabled_doc = "If true, use orbital parameters to compute top of the atmosphere insolation";
    pism_config:surface.debm_simple.paleo.enabled_option = "debm_simple_paleo";
    pism_config:surface.debm_simple.paleo.enabled_type = "flag";

    pism_config:surface.debm_simple.paleo.file = "";
    pism_config:surface.debm_simple.paleo.file_doc = "File containing orbital parameters (:var:`eccentricity`, :var:`obliquity`, :var:`perihelion_longitude`) for paleo-simulations";
    pism_config:surface.debm_simple.paleo.file_option = "debm_simple_paleo_file";
    pism_config:surface.debm_simple.paleo.file_type = "string";

    pism_config:surface.debm_simple.paleo.obliquity =  23.44;
    pism_config:surface.debm_simple.paleo.obliquity_doc = "Mean obliquity (axial tilt) of the Earth";
    pism_config:surface.debm_simple.paleo.obliquity_type = "number";
    pism_config:surface.debm_simple.paleo.obliquity_units = "degree";

    pism_config:surface.debm_simple.paleo.perihelion_longitude =  102.94719;
    pism_config:surface.debm_simple.paleo.perihelion_longitude_doc = "Mean longitude of the perihelion relative to the vernal equinox";
    pism_config:surface.debm_simple.paleo.perihelion_longitude_type = "number";
    pism_config:surface.debm_simple.paleo.perihelion_longitude_units = "degree";

    pism_config:surface.debm_simple.paleo.periodic = "no";
    pism_config:surface.debm_simple.paleo.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.debm_simple.paleo.periodic_type = "flag";

    pism_config:surface.debm_simple.phi =  17.5;
    pism_config:surface.debm_simple.phi_doc = "Threshold solar elevation angle above which melt is possible";
    pism_config:surface.debm_simple.phi_type = "number";
    pism_config:surface.debm_simple.phi_units = "degree";

    pism_config:surface.debm_simple.positive_threshold_temp = 273.15;
    pism_config:surface.debm_simple.positive_threshold_temp_doc = "Temperature threshold used to define the \"positive\" temperature";
    pism_config:surface.debm_simple.positive_threshold_temp_type = "number";
    pism_config:surface.debm_simple.positive_threshold_temp_units = "Kelvin";

    pism_config:surface.debm_simple.refreeze = 0.6;
    pism_config:surface.debm_simple.refreeze_doc = "Refreeze fraction: this fraction of snow melt is assumed to re-freeze. See also :config:`surface.debm_simple.refreeze_ice_melt`.";
    pism_config:surface.debm_simple.refreeze_type = "number";
    pism_config:surface.debm_simple.refreeze_units = "1";

    pism_config:surface.debm_simple.refreeze_ice_melt = "no";
    pism_config:surface.debm_simple.refreeze_ice_melt_doc = "If set to 'yes', refreeze :config:`surface.debm_simple.refreeze` fraction of melted ice, otherwise all of the melted ice runs off.";
    pism_config:surface.debm_simple.refreeze_ice_melt_type = "flag";

    pism_config:surface.debm_simple.solar_constant = 1361.0;
    pism_config:surface.debm_simple.solar_constant_doc = "Mean solar electromagnetic radiation (total solar irradiance) per unit area :cite:`Kopp2011`";
    pism_config:surface.debm_simple.solar_constant_type = "number";
    pism_config:surface.debm_simple.solar_constant_units = "W m-2";

    pism_config:surface.debm_simple.std_dev = 5.0;
    pism_config:surface.debm_simple.std_dev_doc = "Standard deviation of daily near-surface air temperature variation";
    pism_config:surface.debm_simple.std_dev_type = "number";
    pism_config:surface.debm_simple.std_dev_units = "Kelvin";

    pism_config:surface.debm_simple.std_dev.file = "";
    pism_config:surface.debm_simple.std_dev.file_doc = "The file to read :var:`air_temp_sd` (standard deviation of air temperature) from";
    pism_config:surface.debm_simple.std_dev.file_option = "debm_simple_sd_file";
    pism_config:surface.debm_simple.std_dev.file_type = "string";

    pism_config:surface.debm_simple.std_dev.param.a = -0.15;
    pism_config:surface.debm_simple.std_dev.param.a_doc = "Parameter `a` in `\\sigma = \\max(a\\, (T - T_{\\text{melting}}) + b, 0)`. Used only if :config:`surface.debm_simple.std_dev.param.enabled` is set to yes.";
    pism_config:surface.debm_simple.std_dev.param.a_type = "number";
    pism_config:surface.debm_simple.std_dev.param.a_units = "1";

    pism_config:surface.debm_simple.std_dev.param.b = 0.66;
    pism_config:surface.debm_simple.std_dev.param.b_doc = "Parameter `b` in `\\sigma = \\max(a\\, (T - T_{\\text{melting}}) + b, 0)`. Used only if :config:`surface.debm_simple.std_dev.param.enabled` is set to yes.";
    pism_config:surface.debm_simple.std_dev.param.b_type = "number";
    pism_config:surface.debm_simple.std_dev.param.b_units = "Kelvin";

    pism_config:surface.debm_simple.std_dev.param.enabled = "no";
    pism_config:surface.debm_simple.std_dev.param.enabled_doc = "Parameterize standard deviation as a linear function of air temperature over ice-covered grid cells. The region of application is controlled by :config:`geometry.ice_free_thickness_standard`.";
    pism_config:surface.debm_simple.std_dev.param.enabled_type = "flag";

    pism_config:surface.debm_simple.std_dev.periodic = "no";
    pism_config:surface.debm_simple.std_dev.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.debm_simple.std_dev.periodic_type = "flag";

    pism_config:surface.debm_simple.tau_a_intercept = 0.65;
    pism_config:surface.debm_simple.tau_a_intercept_doc = "Intercept in the parametrization of atmosphere transmissivity";
    pism_config:surface.debm_simple.tau_a_intercept_type = "number";
    pism_config:surface.debm_simple.tau_a_intercept_units = "";

    pism_config:surface.debm_simple.tau_a_slope = 0.000032;
    pism_config:surface.debm_simple.tau_a_slope_doc = "Slope in the parametrization of atmosphere transmissivity";
    pism_config:surface.debm_simple.tau_a_slope_type = "number";
    pism_config:surface.debm_simple.tau_a_slope_units = "m-1";

    pism_config:surface.delta_T.file = "";
    pism_config:surface.delta_T.file_doc = "Name of the file containing temperature offsets.";
    pism_config:surface.delta_T.file_option = "surface_delta_T_file";
    pism_config:surface.delta_T.file_type = "string";

    pism_config:surface.delta_T.periodic = "no";
    pism_config:surface.delta_T.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.delta_T.periodic_type = "flag";

    pism_config:surface.elevation_change.file = "";
    pism_config:surface.elevation_change.file_doc = "Name of the file containing the reference surface elevation field (variable :var:`usurf`).";
    pism_config:surface.elevation_change.file_option = "surface_elevation_change_file";
    pism_config:surface.elevation_change.file_type = "string";

    pism_config:surface.elevation_change.periodic = "no";
    pism_config:surface.elevation_change.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.elevation_change.periodic_type = "flag";

    pism_config:surface.elevation_change.smb.exp_factor = 0;
    pism_config:surface.elevation_change.smb.exp_factor_doc = "Exponential for the surface mass balance.";
    pism_config:surface.elevation_change.smb.exp_factor_option = "smb_exp_factor";
    pism_config:surface.elevation_change.smb.exp_factor_type = "number";
    pism_config:surface.elevation_change.smb.exp_factor_units = "Kelvin-1";

    pism_config:surface.elevation_change.smb.lapse_rate = 0;
    pism_config:surface.elevation_change.smb.lapse_rate_doc = "Lapse rate for the surface mass balance.";
    pism_config:surface.elevation_change.smb.lapse_rate_option = "smb_lapse_rate";
    pism_config:surface.elevation_change.smb.lapse_rate_type = "number";
    pism_config:surface.elevation_change.smb.lapse_rate_units = "(m / year) / km";

    pism_config:surface.elevation_change.smb.method = "shift";
    pism_config:surface.elevation_change.smb.method_choices = "scale,shift";
    pism_config:surface.elevation_change.smb.method_doc = "Choose the SMB adjustment method. ``scale``: use temperature-change-dependent scaling factor. ``shift``: use the SMB lapse rate.";
    pism_config:surface.elevation_change.smb.method_option = "smb_adjustment";
    pism_config:surface.elevation_change.smb.method_type = "keyword";

    pism_config:surface.elevation_change.temperature_lapse_rate = 0;
    pism_config:surface.elevation_change.temperature_lapse_rate_doc = "Lapse rate for the temperature at the top of the ice.";
    pism_config:surface.elevation_change.temperature_lapse_rate_option = "temp_lapse_rate";
    pism_config:surface.elevation_change.temperature_lapse_rate_type = "number";
    pism_config:surface.elevation_change.temperature_lapse_rate_units = "K / km";

    pism_config:surface.force_to_thickness.alpha = 0.01;
    pism_config:surface.force_to_thickness.alpha_doc = "exponential coefficient in force-to-thickness mechanism";
    pism_config:surface.force_to_thickness.alpha_option = "force_to_thickness_alpha";
    pism_config:surface.force_to_thickness.alpha_type = "number";
    pism_config:surface.force_to_thickness.alpha_units = "year-1";

    pism_config:surface.force_to_thickness.file = "";
    pism_config:surface.force_to_thickness.file_doc = "The name of the file to read the target ice thickness from.";
    pism_config:surface.force_to_thickness.file_option = "force_to_thickness_file";
    pism_config:surface.force_to_thickness.file_type = "string";

    pism_config:surface.force_to_thickness.ice_free_alpha_factor = 1.0;
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_doc = ":config:`surface.force_to_thickness.alpha` is multiplied by this factor in areas that are ice-free according to the target ice thickness and :config:`surface.force_to_thickness.ice_free_thickness_threshold`";
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_option = "force_to_thickness_ice_free_alpha_factor";
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_type = "number";
    pism_config:surface.force_to_thickness.ice_free_alpha_factor_units = "1";

    pism_config:surface.force_to_thickness.ice_free_thickness_threshold = 1.0;
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_doc = "threshold of ice thickness in the force-to-thickness target field. Used to determine whether to use :config:`surface.force_to_thickness.ice_free_alpha_factor`.";
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_option = "force_to_thickness_ice_free_thickness_threshold";
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_type = "number";
    pism_config:surface.force_to_thickness.ice_free_thickness_threshold_units = "meters";

    pism_config:surface.force_to_thickness.start_time = -4.54e9;
    pism_config:surface.force_to_thickness.start_time_doc = "Starting time for the \"force to thickness\" modifier; the default is \"start from the creation of the Earth.\"";
    pism_config:surface.force_to_thickness.start_time_type = "number";
    pism_config:surface.force_to_thickness.start_time_units = "years";

    pism_config:surface.given.file = "";
    pism_config:surface.given.file_doc = "Name of the file containing climate forcing fields.";
    pism_config:surface.given.file_option = "surface_given_file";
    pism_config:surface.given.file_type = "string";

    pism_config:surface.given.periodic = "no";
    pism_config:surface.given.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.given.periodic_type = "flag";

    pism_config:surface.given.smb_max = 91000;
    pism_config:surface.given.smb_max_doc = "Maximum climatic mass balance value (used to check input data). Corresponds to 100 m/year ice equivalent.";
    pism_config:surface.given.smb_max_type = "number";
    pism_config:surface.given.smb_max_units = "kg m-2 year-1";

    pism_config:surface.ismip6.file = "";
    pism_config:surface.ismip6.file_doc = "Name of the file containing climate forcing anomaly fields.";
    pism_config:surface.ismip6.file_option = "surface_ismip6_file";
    pism_config:surface.ismip6.file_type = "string";

    pism_config:surface.ismip6.periodic = "no";
    pism_config:surface.ismip6.periodic_doc = "If true, interpret forcing data as periodic in time";
    pism_config:surface.ismip6.periodic_type = "flag";

    pism_config:surface.ismip6.reference_file = "";
    pism_config:surface.ismip6.reference_file_doc = "Name of the file containing reference climate forcing fields.";
    pism_config:surface.ismip6.reference_file_option = "surface_ismip6_reference_file";
    pism_config:surface.ismip6.reference_file_type = "string";

    pism_config:surface.mass_balance_year_start_day = 274;
    pism_config:surface.mass_balance_year_start_day_doc = "day of year for October 1st, beginning of the balance year in northern latitudes.";
    pism_config:surface.mass_balance_year_start_day_type = "integer";
    pism_config:surface.mass_balance_year_start_day_units = "ordinal day number";

    pism_config:surface.models = "given";
    pism_config:surface.models_doc = "Comma-separated list of surface models and modifiers";
    pism_config:surface.models_option = "surface";
    pism_config:surface.models_type = "string";

    pism_config:surface.pdd.air_temp_all_precip_as_rain = 275.15;
    pism_config:surface.pdd.air_temp_all_precip_as_rain_doc = "threshold temperature above which all precipitation is rain; must exceed :config:`surface.pdd.air_temp_all_precip_as_snow` to avoid division by zero, because difference is in a denominator";
    pism_config:surface.pdd.air_temp_all_precip_as_rain_type = "number";
    pism_config:surface.pdd.air_temp_all_precip_as_rain_units = "Kelvin";

    pism_config:surface.pdd.air_temp_all_precip_as_snow = 273.15;
    pism_config:surface.pdd.air_temp_all_precip_as_snow_doc = "threshold temperature below which all precipitation is snow";
    pism_config:surface.pdd.air_temp_all_precip_as_snow_type = "number";
    pism_config:surface.pdd.air_temp_all_precip_as_snow_units = "Kelvin";

    pism_config:surface.pdd.factor_ice = 0.00879120879120879;
    pism_config:surface.pdd.factor_ice_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`; = (8 mm liquid-water-equivalent) / (pos degree day)";
    pism_config:surface.pdd.factor_ice_type = "number";
    pism_config:surface.pdd.factor_ice_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.factor_snow = 0.0032967032967033;
    pism_config:surface.pdd.factor_snow_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`; = (3 mm liquid-water-equivalent) / (pos degree day)";
    pism_config:surface.pdd.factor_snow_type = "number";
    pism_config:surface.pdd.factor_snow_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.T_c = 272.15;
    pism_config:surface.pdd.fausto.T_c_doc = "= -1 + 273.15; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.T_c_type = "number";
    pism_config:surface.pdd.fausto.T_c_units = "Kelvin";

    pism_config:surface.pdd.fausto.T_w = 283.15;
    pism_config:surface.pdd.fausto.T_w_doc = "= 10 + 273.15; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.T_w_type = "number";
    pism_config:surface.pdd.fausto.T_w_units = "Kelvin";

    pism_config:surface.pdd.fausto.beta_ice_c = 0.015;
    pism_config:surface.pdd.fausto.beta_ice_c_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.beta_ice_c_type = "number";
    pism_config:surface.pdd.fausto.beta_ice_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_ice_w = 0.007;
    pism_config:surface.pdd.fausto.beta_ice_w_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.beta_ice_w_type = "number";
    pism_config:surface.pdd.fausto.beta_ice_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_snow_c = 0.003;
    pism_config:surface.pdd.fausto.beta_snow_c_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.beta_snow_c_type = "number";
    pism_config:surface.pdd.fausto.beta_snow_c_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.beta_snow_w = 0.003;
    pism_config:surface.pdd.fausto.beta_snow_w_doc = "water-equivalent thickness; for formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.beta_snow_w_type = "number";
    pism_config:surface.pdd.fausto.beta_snow_w_units = "meter / (Kelvin day)";

    pism_config:surface.pdd.fausto.enabled = "false";
    pism_config:surface.pdd.fausto.enabled_doc = "Set PDD parameters using formulas (6) and (7) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.enabled_option = "pdd_fausto";
    pism_config:surface.pdd.fausto.enabled_type = "flag";

    pism_config:surface.pdd.fausto.latitude_beta_w = 72.0;
    pism_config:surface.pdd.fausto.latitude_beta_w_doc = "latitude below which to use warm case, in formula (6) in :cite:`Faustoetal2009`";
    pism_config:surface.pdd.fausto.latitude_beta_w_type = "number";
    pism_config:surface.pdd.fausto.latitude_beta_w_units = "degree_north";

    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio = 0.75;
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_doc = "How much firn as a fraction of accumulation is turned into ice";
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_type = "number";
    pism_config:surface.pdd.firn_compaction_to_accumulation_ratio_units = "1";

    pism_config:surface.pdd.firn_depth_file = "";
    pism_config:surface.pdd.firn_depth_file_doc = "The name of the file to read the firn_depth from.";
    pism_config:surface.pdd.firn_depth_file_option = "pdd_firn_depth_file";
    pism_config:surface.pdd.firn_depth_file_type = "string";

    pism_config:surface.pdd.interpret_precip_as_snow = "no";
    pism_config:surface.pdd.interpret_precip_as_snow_doc = "Interpret precipitation as snow fall.";
    pism_config:surface.pdd.interpret_precip_as_snow_type = "flag";

    pism_config:surface.pdd.max_evals_per_year = 52;
    pism_config:surface.pdd.max_evals_per_year_doc = "maximum number of times the PDD scheme will ask for air temperature and precipitation to build location-dependent time series for computing (expected) number of positive degree days and snow accumulation; the default means the PDD uses weekly samples of the annual cycle; see also :config:`surface.pdd.std_dev.value`";
    pism_config:surface.pdd.max_evals_per_year_type = "integer";
    pism_config:surface.pdd.max_evals_per_year_units = "count";

    pism_config:surface.pdd.method = "expectation_integral";
    pism_config:surface.pdd.method_choices = "expectation_integral,repeatable_random_process,random_process";
    pism_config:surface.pdd.method_doc = "PDD implementation method";
    pism_config:surface.pdd.method_option = "pdd_method";
    pism_config:surface.pdd.method_type = "keyword";

    pism_config:surface.pdd.positive_threshold_temp = 273.15;
    pism_config:surface.pdd.positive_threshold_temp_doc = "temperature used to determine meaning of \"positive\" degree day";
    pism_config:surface.pdd.positive_threshold_temp_type = "number";
    pism_config:surface.pdd.positive_threshold_temp_units = "Kelvin";

    pism_config:surface.pdd.refreeze = 0.6;
    pism_config:surface.pdd.refreeze_doc = "EISMINT-Greenland value :cite:`RitzEISMINT`";
    pism_config:surface.pdd.refreeze_type = "number";
    pism_config:surface.pdd.refreeze_units = "1";

    pism_config:surface.pdd.refreeze_ice_melt = "yes";
    pism_config:surface.pdd.refreeze_ice_melt_doc = "If set to \"yes\", refreeze :config:`surface.pdd.refreeze` fraction of melted ice, otherwise all of the melted ice runs off.";
    pism_config:surface.pdd.refreeze_ice_melt_type = "flag";

    pism_config:surface.pdd.std_dev.file = "";
    pism_config:surface.pdd.std_dev.file_doc = "The name of the file to read ``air_temp_sd`` (standard deviation of air temperature) from.";
    pism_config:surface.pdd.std_dev.file_option = "pdd_sd_file";
    pism_config:surface.pdd.std_dev.file_type = "string";

    pism_config:surface.pdd.std_dev.lapse_lat_base = 72.0;
    pism_config:surface.pdd.std_dev.lapse_lat_base_doc = "standard deviationis is a function of latitude, with value :config:`surface.pdd.std_dev.value` at this latitude; this value is only active if :config:`surface.pdd.std_dev.lapse_lat_rate` is nonzero";
    pism_config:surface.pdd.std_dev.lapse_lat_base_type = "number";
    pism_config:surface.pdd.std_dev.lapse_lat_base_units = "degree_north";

    pism_config:surface.pdd.std_dev.lapse_lat_rate = 0.0;
    pism_config:surface.pdd.std_dev.lapse_lat_rate_doc = "standard deviation is a function of latitude, with rate of change with respect to latitude given by this constant";
    pism_config:surface.pdd.std_dev.lapse_lat_rate_type = "number";
    pism_config:surface.pdd.std_dev.lapse_lat_rate_units = "Kelvin / degree_north";

    pism_config:surface.pdd.std_dev.param_a = -0.15;
    pism_config:surface.pdd.std_dev.param_a_doc = "Parameter `a` in `\\Sigma = aT + b`, with `T` in degrees C. Used only if :config:`surface.pdd.std_dev.use_param` is set to yes.";
    pism_config:surface.pdd.std_dev.param_a_type = "number";
    pism_config:surface.pdd.std_dev.param_a_units = "pure number";

    pism_config:surface.pdd.std_dev.param_b = 0.66;
    pism_config:surface.pdd.std_dev.param_b_doc = "Parameter `b` in `\\Sigma = aT + b`, with `T` in degrees C. Used only if :config:`surface.pdd.std_dev.use_param` is set to yes.";
    pism_config:surface.pdd.std_dev.param_b_type = "number";
    pism_config:surface.pdd.std_dev.param_b_units = "Kelvin";

    pism_config:surface.pdd.std_dev.periodic = "no";
    pism_config:surface.pdd.std_dev.periodic_doc = "If true, interpret ``air_temp_sd`` read from :config:`surface.pdd.std_dev.file` as periodic in time";
    pism_config:surface.pdd.std_dev.periodic_type = "flag";

    pism_config:surface.pdd.std_dev.use_param = "no";
    pism_config:surface.pdd.std_dev.use_param_doc = "Parameterize standard deviation as a linear function of air temperature over ice-covered grid cells. The region of application is controlled by :config:`geometry.ice_free_thickness_standard`.";
    pism_config:surface.pdd.std_dev.use_param_type = "flag";

    pism_config:surface.pdd.std_dev.value = 5.0;
    pism_config:surface.pdd.std_dev.value_doc = "standard deviation of daily temp variation; = EISMINT-Greenland value :cite:`RitzEISMINT`";
    pism_config:surface.pdd.std_dev.value_type = "number";
    pism_config:surface.pdd.std_dev.value_units = "Kelvin";

    pism_config:surface.pressure = 0.0;
    pism_config:surface.pressure_doc = "atmospheric pressure; = pressure at ice surface";
    pism_config:surface.pressure_type = "number";
    pism_config:surface.pressure_units = "Pascal";

    pism_config:surface.temp_to_runoff_a = 0.5;
    pism_config:surface.temp_to_runoff_a_doc = "a in runoff=a * temp + b";
    pism_config:surface.temp_to_runoff_a_type = "number";
    pism_config:surface.temp_to_runoff_a_units = "K-1";

    pism_config:time.calendar = "365_day";
    pism_config:time.calendar_choices = "standard,gregorian,proleptic_gregorian,noleap,365_day,360_day,julian";
    pism_config:time.calendar_doc = "The calendar to use.";
    pism_config:time.calendar_option = "calendar";
    pism_config:time.calendar_type = "keyword";

    pism_config:time.dimension_name = "time";
    pism_config:time.dimension_name_doc = "The name of the time dimension in PISM output files.";
    pism_config:time.dimension_name_type = "string";

    pism_config:time.eemian_end = -114500.0;
    pism_config:time.eemian_end_doc = "End of the Eemian interglacial period. See :cite:`Greve97Greenland`.";
    pism_config:time.eemian_end_type = "number";
    pism_config:time.eemian_end_units = "years";

    pism_config:time.eemian_start = -132000.0;
    pism_config:time.eemian_start_doc = "Start of the Eemian interglacial period. See :cite:`Greve97Greenland`.";
    pism_config:time.eemian_start_type = "number";
    pism_config:time.eemian_start_units = "years";

    pism_config:time.end = "";
    pism_config:time.end_doc = "End time, interpreted relative to :config:`time.reference_date`.";
    pism_config:time.end_option = "ye";
    pism_config:time.end_type = "string";

    pism_config:time.file = "";
    pism_config:time.file_doc = "Name of the file used to set :config:`time.start`, :config:`time.end`, :config:`time.calendar`, and :config:`time.reference_date`";
    pism_config:time.file_type = "string";
    pism_config:time.file_option = "time_file";

    pism_config:time.file.continue = "false";
    pism_config:time.file.continue_doc = "If true, don't set :config:`time.start` using :config:`time.file` (helpful when continuing an interrupted simulation)";
    pism_config:time.file.continue_type = "flag";

    pism_config:time.holocene_start = -11000.0;
    pism_config:time.holocene_start_doc = "Start of the Holocene interglacial period. See :cite:`Greve97Greenland`.";
    pism_config:time.holocene_start_type = "number";
    pism_config:time.holocene_start_units = "years";

    pism_config:time.reference_date = "0001-1-1";
    pism_config:time.reference_date_doc = "year-month-day; reference date used for calendar computations and in PISM output files";
    pism_config:time.reference_date_type = "string";

    pism_config:time.run_length = 1000;
    pism_config:time.run_length_doc = "Run length";
    pism_config:time.run_length_option = "y";
    pism_config:time.run_length_type = "number";
    pism_config:time.run_length_units = "365days";

    pism_config:time.start = "";
    pism_config:time.start_doc = "Start time, interpreted relative to :config:`time.reference_date`.";
    pism_config:time.start_option = "ys";
    pism_config:time.start_type = "string";

    pism_config:time_stepping.adaptive_ratio = 0.12;
    pism_config:time_stepping.adaptive_ratio_doc = "Adaptive time stepping ratio for the explicit scheme for the mass balance equation; :cite:`BBL`, inequality (25)";
    pism_config:time_stepping.adaptive_ratio_option = "adapt_ratio";
    pism_config:time_stepping.adaptive_ratio_type = "number";
    pism_config:time_stepping.adaptive_ratio_units = "1";

    pism_config:time_stepping.assume_bed_elevation_changed = "no";
    pism_config:time_stepping.assume_bed_elevation_changed_doc = "If set, assume that bed elevation changes every time step. If not set, PISM tries to avoid unnecessary computations if the bed deformation model did not update bed elevation (to reduce the computational cost a little bit).";
    pism_config:time_stepping.assume_bed_elevation_changed_type = "flag";

    pism_config:time_stepping.hit_extra_times = "yes";
    pism_config:time_stepping.hit_extra_times_doc = "Modify the time-stepping mechanism to hit times requested using :config:`output.extra.times`.";
    pism_config:time_stepping.hit_extra_times_option = "extra_force_output_times";
    pism_config:time_stepping.hit_extra_times_type = "flag";

    pism_config:time_stepping.hit_multiples = 0.0;
    pism_config:time_stepping.hit_multiples_doc = "Hit every X years, where X is specified using this parameter. Use 0 to disable.";
    pism_config:time_stepping.hit_multiples_option = "timestep_hit_multiples";
    pism_config:time_stepping.hit_multiples_type = "integer";
    pism_config:time_stepping.hit_multiples_units = "years";

    pism_config:time_stepping.hit_save_times = "no";
    pism_config:time_stepping.hit_save_times_doc = "Modify the time-stepping mechanism to hit times requested using :config:`output.snapshot.times`.";
    pism_config:time_stepping.hit_save_times_option = "save_force_output_times";
    pism_config:time_stepping.hit_save_times_type = "flag";

    pism_config:time_stepping.hit_ts_times = "no";
    pism_config:time_stepping.hit_ts_times_doc = "Modify the time-stepping mechanism to hit times requested using :config:`output.timeseries.times`.";
    pism_config:time_stepping.hit_ts_times_type = "flag";

    pism_config:time_stepping.maximum_time_step = 60.0;
    pism_config:time_stepping.maximum_time_step_doc = "Maximum allowed time step length";
    pism_config:time_stepping.maximum_time_step_option = "max_dt";
    pism_config:time_stepping.maximum_time_step_type = "number";
    pism_config:time_stepping.maximum_time_step_units = "365days";

    pism_config:time_stepping.resolution = 1.0;
    pism_config:time_stepping.resolution_doc = "Time steps are rounded down to be a multiple of this number (set to zero to allow arbitrary time step lengths)";
    pism_config:time_stepping.resolution_type = "number";
    pism_config:time_stepping.resolution_units = "seconds";

    pism_config:time_stepping.skip.enabled = "no";
    pism_config:time_stepping.skip.enabled_doc = "Use the temperature, age, and SSA stress balance computation skipping mechanism.";
    pism_config:time_stepping.skip.enabled_option = "skip";
    pism_config:time_stepping.skip.enabled_type = "flag";

    pism_config:time_stepping.skip.max = 10;
    pism_config:time_stepping.skip.max_doc = "Number of mass-balance steps, including SIA diffusivity updates, to perform before a the temperature, age, and SSA stress balance computations are done";
    pism_config:time_stepping.skip.max_option = "skip_max";
    pism_config:time_stepping.skip.max_type = "integer";
    pism_config:time_stepping.skip.max_units = "count";

    pism_config:long_name = "PISM configuration flags and parameters.";
    pism_config:long_name_doc = "The long_name attribute is required by CF conventions. It is not used by PISM itself.";
}
