netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:ocean_kill  = "true";
    pism_overrides:ocean_kill_doc = "If used with input from a NetCDF initialization file which has ice-free ocean mask, will zero out ice thicknesses in areas that were ice-free ocean at time zero. This is calving at the location of the original calving front.";

    pism_overrides:bootstrapping_geothermal_flux_value_no_var = 0.050;
    pism_overrides:bootstrapping_geothermal_flux_value_no_var_doc = "W m-2; geothermal flux value to use if bheatflx variable is absent in bootstrapping file";

    pism_overrides:pdd_std_dev = 5.0;
    pism_overrides:pdd_std_dev_doc = "K; std dev of daily temp variation; value from [\\ref RitzEISMINT] ";


   pism_overrides:institution = "University of Alaska Fairbanks";
   pism_overrides:institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";

    pism_overrides:enhancement_factor = 3.0;
    pism_overrides:enhancement_factor_doc = "; Flow enhancement factor for SIA";

}
